module DotProductModule_1(input clk,
    input [17:0] io_a_11,
    input [17:0] io_a_10,
    input [17:0] io_a_9,
    input [17:0] io_a_8,
    input [17:0] io_a_7,
    input [17:0] io_a_6,
    input [17:0] io_a_5,
    input [17:0] io_a_4,
    input [17:0] io_a_3,
    input [17:0] io_a_2,
    input [17:0] io_a_1,
    input [17:0] io_a_0,
    input [17:0] io_b_11,
    input [17:0] io_b_10,
    input [17:0] io_b_9,
    input [17:0] io_b_8,
    input [17:0] io_b_7,
    input [17:0] io_b_6,
    input [17:0] io_b_5,
    input [17:0] io_b_4,
    input [17:0] io_b_3,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    output[17:0] io_o
);

  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  wire[17:0] T3;
  wire[17:0] T4;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  wire[17:0] T8;
  reg [17:0] R9;
  wire[17:0] T10;
  wire[17:0] T116;
  wire[21:0] T11;
  wire[35:0] T12;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  reg [17:0] R16;
  wire[17:0] T17;
  wire[17:0] T117;
  wire[21:0] T18;
  wire[35:0] T19;
  wire[17:0] T20;
  wire[17:0] T21;
  wire[17:0] T22;
  wire[17:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;
  reg [17:0] R26;
  wire[17:0] T27;
  wire[17:0] T118;
  wire[21:0] T28;
  wire[35:0] T29;
  wire[17:0] T30;
  wire[17:0] T31;
  wire[17:0] T32;
  reg [17:0] R33;
  wire[17:0] T34;
  wire[17:0] T119;
  wire[21:0] T35;
  wire[35:0] T36;
  wire[17:0] T37;
  wire[17:0] T38;
  wire[17:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  wire[17:0] T42;
  wire[17:0] T43;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[17:0] T46;
  wire[17:0] T47;
  wire[17:0] T48;
  reg [17:0] R49;
  wire[17:0] T50;
  wire[17:0] T120;
  wire[21:0] T51;
  wire[35:0] T52;
  wire[17:0] T53;
  wire[17:0] T54;
  wire[17:0] T55;
  reg [17:0] R56;
  wire[17:0] T57;
  wire[17:0] T121;
  wire[21:0] T58;
  wire[35:0] T59;
  wire[17:0] T60;
  wire[17:0] T61;
  wire[17:0] T62;
  wire[17:0] T63;
  wire[17:0] T64;
  wire[17:0] T65;
  reg [17:0] R66;
  wire[17:0] T67;
  wire[17:0] T122;
  wire[21:0] T68;
  wire[35:0] T69;
  wire[17:0] T70;
  wire[17:0] T71;
  wire[17:0] T72;
  reg [17:0] R73;
  wire[17:0] T74;
  wire[17:0] T123;
  wire[21:0] T75;
  wire[35:0] T76;
  wire[17:0] T77;
  wire[17:0] T78;
  wire[17:0] T79;
  wire[17:0] T80;
  wire[17:0] T81;
  wire[17:0] T82;
  wire[17:0] T83;
  wire[17:0] T84;
  wire[17:0] T85;
  reg [17:0] R86;
  wire[17:0] T87;
  wire[17:0] T124;
  wire[21:0] T88;
  wire[35:0] T89;
  wire[17:0] T90;
  wire[17:0] T91;
  wire[17:0] T92;
  reg [17:0] R93;
  wire[17:0] T94;
  wire[17:0] T125;
  wire[21:0] T95;
  wire[35:0] T96;
  wire[17:0] T97;
  wire[17:0] T98;
  wire[17:0] T99;
  wire[17:0] T100;
  wire[17:0] T101;
  wire[17:0] T102;
  reg [17:0] R103;
  wire[17:0] T104;
  wire[17:0] T126;
  wire[21:0] T105;
  wire[35:0] T106;
  wire[17:0] T107;
  wire[17:0] T108;
  wire[17:0] T109;
  reg [17:0] R110;
  wire[17:0] T111;
  wire[17:0] T127;
  wire[21:0] T112;
  wire[35:0] T113;
  wire[17:0] T114;
  wire[17:0] T115;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R9 = {1{$random}};
    R16 = {1{$random}};
    R26 = {1{$random}};
    R33 = {1{$random}};
    R49 = {1{$random}};
    R56 = {1{$random}};
    R66 = {1{$random}};
    R73 = {1{$random}};
    R86 = {1{$random}};
    R93 = {1{$random}};
    R103 = {1{$random}};
    R110 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_o = T0;
  assign T0 = T1;
  assign T1 = T39 + T2;
  assign T2 = T3;
  assign T3 = T4;
  assign T4 = T22 + T5;
  assign T5 = T6;
  assign T6 = T7;
  assign T7 = T15 + T8;
  assign T8 = R9;
  assign T10 = T116;
  assign T116 = T11[5'h11:1'h0];
  assign T11 = $signed(T12) >>> 4'he;
  assign T12 = $signed(T14) * $signed(T13);
  assign T13 = io_b_11;
  assign T14 = io_a_11;
  assign T15 = R16;
  assign T17 = T117;
  assign T117 = T18[5'h11:1'h0];
  assign T18 = $signed(T19) >>> 4'he;
  assign T19 = $signed(T21) * $signed(T20);
  assign T20 = io_b_10;
  assign T21 = io_a_10;
  assign T22 = T23;
  assign T23 = T24;
  assign T24 = T32 + T25;
  assign T25 = R26;
  assign T27 = T118;
  assign T118 = T28[5'h11:1'h0];
  assign T28 = $signed(T29) >>> 4'he;
  assign T29 = $signed(T31) * $signed(T30);
  assign T30 = io_b_9;
  assign T31 = io_a_9;
  assign T32 = R33;
  assign T34 = T119;
  assign T119 = T35[5'h11:1'h0];
  assign T35 = $signed(T36) >>> 4'he;
  assign T36 = $signed(T38) * $signed(T37);
  assign T37 = io_b_8;
  assign T38 = io_a_8;
  assign T39 = T40;
  assign T40 = T41;
  assign T41 = T79 + T42;
  assign T42 = T43;
  assign T43 = T44;
  assign T44 = T62 + T45;
  assign T45 = T46;
  assign T46 = T47;
  assign T47 = T55 + T48;
  assign T48 = R49;
  assign T50 = T120;
  assign T120 = T51[5'h11:1'h0];
  assign T51 = $signed(T52) >>> 4'he;
  assign T52 = $signed(T54) * $signed(T53);
  assign T53 = io_b_7;
  assign T54 = io_a_7;
  assign T55 = R56;
  assign T57 = T121;
  assign T121 = T58[5'h11:1'h0];
  assign T58 = $signed(T59) >>> 4'he;
  assign T59 = $signed(T61) * $signed(T60);
  assign T60 = io_b_6;
  assign T61 = io_a_6;
  assign T62 = T63;
  assign T63 = T64;
  assign T64 = T72 + T65;
  assign T65 = R66;
  assign T67 = T122;
  assign T122 = T68[5'h11:1'h0];
  assign T68 = $signed(T69) >>> 4'he;
  assign T69 = $signed(T71) * $signed(T70);
  assign T70 = io_b_5;
  assign T71 = io_a_5;
  assign T72 = R73;
  assign T74 = T123;
  assign T123 = T75[5'h11:1'h0];
  assign T75 = $signed(T76) >>> 4'he;
  assign T76 = $signed(T78) * $signed(T77);
  assign T77 = io_b_4;
  assign T78 = io_a_4;
  assign T79 = T80;
  assign T80 = T81;
  assign T81 = T99 + T82;
  assign T82 = T83;
  assign T83 = T84;
  assign T84 = T92 + T85;
  assign T85 = R86;
  assign T87 = T124;
  assign T124 = T88[5'h11:1'h0];
  assign T88 = $signed(T89) >>> 4'he;
  assign T89 = $signed(T91) * $signed(T90);
  assign T90 = io_b_3;
  assign T91 = io_a_3;
  assign T92 = R93;
  assign T94 = T125;
  assign T125 = T95[5'h11:1'h0];
  assign T95 = $signed(T96) >>> 4'he;
  assign T96 = $signed(T98) * $signed(T97);
  assign T97 = io_b_2;
  assign T98 = io_a_2;
  assign T99 = T100;
  assign T100 = T101;
  assign T101 = T109 + T102;
  assign T102 = R103;
  assign T104 = T126;
  assign T126 = T105[5'h11:1'h0];
  assign T105 = $signed(T106) >>> 4'he;
  assign T106 = $signed(T108) * $signed(T107);
  assign T107 = io_b_1;
  assign T108 = io_a_1;
  assign T109 = R110;
  assign T111 = T127;
  assign T127 = T112[5'h11:1'h0];
  assign T112 = $signed(T113) >>> 4'he;
  assign T113 = $signed(T115) * $signed(T114);
  assign T114 = io_b_0;
  assign T115 = io_a_0;

  always @(posedge clk) begin
    R9 <= T10;
    R16 <= T17;
    R26 <= T27;
    R33 <= T34;
    R49 <= T50;
    R56 <= T57;
    R66 <= T67;
    R73 <= T74;
    R86 <= T87;
    R93 <= T94;
    R103 <= T104;
    R110 <= T111;
  end
endmodule

module MatrixVectorMultModule_1(input clk,
    input [17:0] io_a_2_11,
    input [17:0] io_a_2_10,
    input [17:0] io_a_2_9,
    input [17:0] io_a_2_8,
    input [17:0] io_a_2_7,
    input [17:0] io_a_2_6,
    input [17:0] io_a_2_5,
    input [17:0] io_a_2_4,
    input [17:0] io_a_2_3,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_11,
    input [17:0] io_a_1_10,
    input [17:0] io_a_1_9,
    input [17:0] io_a_1_8,
    input [17:0] io_a_1_7,
    input [17:0] io_a_1_6,
    input [17:0] io_a_1_5,
    input [17:0] io_a_1_4,
    input [17:0] io_a_1_3,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_11,
    input [17:0] io_a_0_10,
    input [17:0] io_a_0_9,
    input [17:0] io_a_0_8,
    input [17:0] io_a_0_7,
    input [17:0] io_a_0_6,
    input [17:0] io_a_0_5,
    input [17:0] io_a_0_4,
    input [17:0] io_a_0_3,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_b_11,
    input [17:0] io_b_10,
    input [17:0] io_b_9,
    input [17:0] io_b_8,
    input [17:0] io_b_7,
    input [17:0] io_b_6,
    input [17:0] io_b_5,
    input [17:0] io_b_4,
    input [17:0] io_b_3,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] R0;
  reg [17:0] R1;
  reg [17:0] R2;
  wire[17:0] DotProductModule_io_o;
  wire[17:0] DotProductModule_1_io_o;
  wire[17:0] DotProductModule_2_io_o;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
    R2 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_o_0 = R0;
  assign io_o_1 = R1;
  assign io_o_2 = R2;
  DotProductModule_1 DotProductModule(.clk(clk),
       .io_a_11( io_a_0_11 ),
       .io_a_10( io_a_0_10 ),
       .io_a_9( io_a_0_9 ),
       .io_a_8( io_a_0_8 ),
       .io_a_7( io_a_0_7 ),
       .io_a_6( io_a_0_6 ),
       .io_a_5( io_a_0_5 ),
       .io_a_4( io_a_0_4 ),
       .io_a_3( io_a_0_3 ),
       .io_a_2( io_a_0_2 ),
       .io_a_1( io_a_0_1 ),
       .io_a_0( io_a_0_0 ),
       .io_b_11( io_b_11 ),
       .io_b_10( io_b_10 ),
       .io_b_9( io_b_9 ),
       .io_b_8( io_b_8 ),
       .io_b_7( io_b_7 ),
       .io_b_6( io_b_6 ),
       .io_b_5( io_b_5 ),
       .io_b_4( io_b_4 ),
       .io_b_3( io_b_3 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_io_o )
  );
  DotProductModule_1 DotProductModule_1(.clk(clk),
       .io_a_11( io_a_1_11 ),
       .io_a_10( io_a_1_10 ),
       .io_a_9( io_a_1_9 ),
       .io_a_8( io_a_1_8 ),
       .io_a_7( io_a_1_7 ),
       .io_a_6( io_a_1_6 ),
       .io_a_5( io_a_1_5 ),
       .io_a_4( io_a_1_4 ),
       .io_a_3( io_a_1_3 ),
       .io_a_2( io_a_1_2 ),
       .io_a_1( io_a_1_1 ),
       .io_a_0( io_a_1_0 ),
       .io_b_11( io_b_11 ),
       .io_b_10( io_b_10 ),
       .io_b_9( io_b_9 ),
       .io_b_8( io_b_8 ),
       .io_b_7( io_b_7 ),
       .io_b_6( io_b_6 ),
       .io_b_5( io_b_5 ),
       .io_b_4( io_b_4 ),
       .io_b_3( io_b_3 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_1_io_o )
  );
  DotProductModule_1 DotProductModule_2(.clk(clk),
       .io_a_11( io_a_2_11 ),
       .io_a_10( io_a_2_10 ),
       .io_a_9( io_a_2_9 ),
       .io_a_8( io_a_2_8 ),
       .io_a_7( io_a_2_7 ),
       .io_a_6( io_a_2_6 ),
       .io_a_5( io_a_2_5 ),
       .io_a_4( io_a_2_4 ),
       .io_a_3( io_a_2_3 ),
       .io_a_2( io_a_2_2 ),
       .io_a_1( io_a_2_1 ),
       .io_a_0( io_a_2_0 ),
       .io_b_11( io_b_11 ),
       .io_b_10( io_b_10 ),
       .io_b_9( io_b_9 ),
       .io_b_8( io_b_8 ),
       .io_b_7( io_b_7 ),
       .io_b_6( io_b_6 ),
       .io_b_5( io_b_5 ),
       .io_b_4( io_b_4 ),
       .io_b_3( io_b_3 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_2_io_o )
  );

  always @(posedge clk) begin
    R0 <= DotProductModule_io_o;
    R1 <= DotProductModule_1_io_o;
    R2 <= DotProductModule_2_io_o;
  end
endmodule

module DotProductModule_0(input clk,
    input [17:0] io_a_2,
    input [17:0] io_a_1,
    input [17:0] io_a_0,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    output[17:0] io_o
);

  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  reg [17:0] R3;
  wire[17:0] T4;
  wire[17:0] T26;
  wire[21:0] T5;
  wire[35:0] T6;
  wire[17:0] T7;
  wire[17:0] T8;
  wire[17:0] T9;
  wire[17:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  reg [17:0] R13;
  wire[17:0] T14;
  wire[17:0] T27;
  wire[21:0] T15;
  wire[35:0] T16;
  wire[17:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  reg [17:0] R20;
  wire[17:0] T21;
  wire[17:0] T28;
  wire[21:0] T22;
  wire[35:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R3 = {1{$random}};
    R13 = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_o = T0;
  assign T0 = T1;
  assign T1 = T9 + T2;
  assign T2 = R3;
  assign T4 = T26;
  assign T26 = T5[5'h11:1'h0];
  assign T5 = $signed(T6) >>> 4'he;
  assign T6 = $signed(T8) * $signed(T7);
  assign T7 = io_b_2;
  assign T8 = io_a_2;
  assign T9 = T10;
  assign T10 = T11;
  assign T11 = T19 + T12;
  assign T12 = R13;
  assign T14 = T27;
  assign T27 = T15[5'h11:1'h0];
  assign T15 = $signed(T16) >>> 4'he;
  assign T16 = $signed(T18) * $signed(T17);
  assign T17 = io_b_1;
  assign T18 = io_a_1;
  assign T19 = R20;
  assign T21 = T28;
  assign T28 = T22[5'h11:1'h0];
  assign T22 = $signed(T23) >>> 4'he;
  assign T23 = $signed(T25) * $signed(T24);
  assign T24 = io_b_0;
  assign T25 = io_a_0;

  always @(posedge clk) begin
    R3 <= T4;
    R13 <= T14;
    R20 <= T21;
  end
endmodule

module MatrixVectorMultModule_0(input clk,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] R0;
  reg [17:0] R1;
  reg [17:0] R2;
  wire[17:0] DotProductModule_io_o;
  wire[17:0] DotProductModule_1_io_o;
  wire[17:0] DotProductModule_2_io_o;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
    R2 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_o_0 = R0;
  assign io_o_1 = R1;
  assign io_o_2 = R2;
  DotProductModule_0 DotProductModule(.clk(clk),
       .io_a_2( io_a_0_2 ),
       .io_a_1( io_a_0_1 ),
       .io_a_0( io_a_0_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_io_o )
  );
  DotProductModule_0 DotProductModule_1(.clk(clk),
       .io_a_2( io_a_1_2 ),
       .io_a_1( io_a_1_1 ),
       .io_a_0( io_a_1_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_1_io_o )
  );
  DotProductModule_0 DotProductModule_2(.clk(clk),
       .io_a_2( io_a_2_2 ),
       .io_a_1( io_a_2_1 ),
       .io_a_0( io_a_2_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_2_io_o )
  );

  always @(posedge clk) begin
    R0 <= DotProductModule_io_o;
    R1 <= DotProductModule_1_io_o;
    R2 <= DotProductModule_2_io_o;
  end
endmodule

module gModule(
    input [17:0] io_in,
    input [17:0] io_hi,
    input [17:0] io_lo,
    output[17:0] io_ou
);

  wire[17:0] T0;
  wire[17:0] T1;
  wire T2;
  wire[17:0] T3;
  wire[17:0] T4;
  wire T5;
  wire[17:0] T6;
  wire[17:0] T7;


  assign io_ou = T0;
  assign T0 = T5 ? io_hi : T1;
  assign T1 = T2 ? io_lo : io_in;
  assign T2 = $signed(T4) < $signed(T3);
  assign T3 = io_lo;
  assign T4 = io_in;
  assign T5 = $signed(T7) < $signed(T6);
  assign T6 = io_in;
  assign T7 = io_hi;
endmodule

module XNetModule(input clk,
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_y_11,
    input [17:0] io_y_10,
    input [17:0] io_y_9,
    input [17:0] io_y_8,
    input [17:0] io_y_7,
    input [17:0] io_y_6,
    input [17:0] io_y_5,
    input [17:0] io_y_4,
    input [17:0] io_y_3,
    input [17:0] io_y_2,
    input [17:0] io_y_1,
    input [17:0] io_y_0,
    input [17:0] io_z_2,
    input [17:0] io_z_1,
    input [17:0] io_z_0,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_c_2_2,
    input [17:0] io_c_2_1,
    input [17:0] io_c_2_0,
    input [17:0] io_c_1_2,
    input [17:0] io_c_1_1,
    input [17:0] io_c_1_0,
    input [17:0] io_c_0_2,
    input [17:0] io_c_0_1,
    input [17:0] io_c_0_0,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] x_stage_2;
  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  reg [17:0] cz_2;
  wire[17:0] T3;
  reg [17:0] xay_2;
  wire[17:0] T4;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  reg [17:0] x_delay_2;
  reg [17:0] R8;
  reg [17:0] x_stage_1;
  wire[17:0] T9;
  wire[17:0] T10;
  wire[17:0] T11;
  reg [17:0] cz_1;
  wire[17:0] T12;
  reg [17:0] xay_1;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  wire[17:0] T16;
  reg [17:0] x_delay_1;
  reg [17:0] R17;
  reg [17:0] x_stage_0;
  wire[17:0] T18;
  wire[17:0] T19;
  wire[17:0] T20;
  reg [17:0] cz_0;
  wire[17:0] T21;
  reg [17:0] xay_0;
  wire[17:0] T22;
  wire[17:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;
  reg [17:0] x_delay_0;
  reg [17:0] R26;
  wire[17:0] gModule_io_ou;
  wire[17:0] gModule_1_io_ou;
  wire[17:0] gModule_2_io_ou;
  wire[17:0] MatrixVectorMultModule_io_o_2;
  wire[17:0] MatrixVectorMultModule_io_o_1;
  wire[17:0] MatrixVectorMultModule_io_o_0;
  wire[17:0] MatrixVectorMultModule_1_io_o_2;
  wire[17:0] MatrixVectorMultModule_1_io_o_1;
  wire[17:0] MatrixVectorMultModule_1_io_o_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    x_stage_2 = {1{$random}};
    cz_2 = {1{$random}};
    xay_2 = {1{$random}};
    x_delay_2 = {1{$random}};
    R8 = {1{$random}};
    x_stage_1 = {1{$random}};
    cz_1 = {1{$random}};
    xay_1 = {1{$random}};
    x_delay_1 = {1{$random}};
    R17 = {1{$random}};
    x_stage_0 = {1{$random}};
    cz_0 = {1{$random}};
    xay_0 = {1{$random}};
    x_delay_0 = {1{$random}};
    R26 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T1;
  assign T1 = T3 + T2;
  assign T2 = cz_2;
  assign T3 = xay_2;
  assign T4 = T5;
  assign T5 = T7 - T6;
  assign T6 = MatrixVectorMultModule_io_o_2;
  assign T7 = x_delay_2;
  assign T9 = T10;
  assign T10 = T12 + T11;
  assign T11 = cz_1;
  assign T12 = xay_1;
  assign T13 = T14;
  assign T14 = T16 - T15;
  assign T15 = MatrixVectorMultModule_io_o_1;
  assign T16 = x_delay_1;
  assign T18 = T19;
  assign T19 = T21 + T20;
  assign T20 = cz_0;
  assign T21 = xay_0;
  assign T22 = T23;
  assign T23 = T25 - T24;
  assign T24 = MatrixVectorMultModule_io_o_0;
  assign T25 = x_delay_0;
  assign io_o_0 = gModule_io_ou;
  assign io_o_1 = gModule_1_io_ou;
  assign io_o_2 = gModule_2_io_ou;
  MatrixVectorMultModule_1 MatrixVectorMultModule(.clk(clk),
       .io_a_2_11( io_a_11_2 ),
       .io_a_2_10( io_a_10_2 ),
       .io_a_2_9( io_a_9_2 ),
       .io_a_2_8( io_a_8_2 ),
       .io_a_2_7( io_a_7_2 ),
       .io_a_2_6( io_a_6_2 ),
       .io_a_2_5( io_a_5_2 ),
       .io_a_2_4( io_a_4_2 ),
       .io_a_2_3( io_a_3_2 ),
       .io_a_2_2( io_a_2_2 ),
       .io_a_2_1( io_a_1_2 ),
       .io_a_2_0( io_a_0_2 ),
       .io_a_1_11( io_a_11_1 ),
       .io_a_1_10( io_a_10_1 ),
       .io_a_1_9( io_a_9_1 ),
       .io_a_1_8( io_a_8_1 ),
       .io_a_1_7( io_a_7_1 ),
       .io_a_1_6( io_a_6_1 ),
       .io_a_1_5( io_a_5_1 ),
       .io_a_1_4( io_a_4_1 ),
       .io_a_1_3( io_a_3_1 ),
       .io_a_1_2( io_a_2_1 ),
       .io_a_1_1( io_a_1_1 ),
       .io_a_1_0( io_a_0_1 ),
       .io_a_0_11( io_a_11_0 ),
       .io_a_0_10( io_a_10_0 ),
       .io_a_0_9( io_a_9_0 ),
       .io_a_0_8( io_a_8_0 ),
       .io_a_0_7( io_a_7_0 ),
       .io_a_0_6( io_a_6_0 ),
       .io_a_0_5( io_a_5_0 ),
       .io_a_0_4( io_a_4_0 ),
       .io_a_0_3( io_a_3_0 ),
       .io_a_0_2( io_a_2_0 ),
       .io_a_0_1( io_a_1_0 ),
       .io_a_0_0( io_a_0_0 ),
       .io_b_11( io_y_11 ),
       .io_b_10( io_y_10 ),
       .io_b_9( io_y_9 ),
       .io_b_8( io_y_8 ),
       .io_b_7( io_y_7 ),
       .io_b_6( io_y_6 ),
       .io_b_5( io_y_5 ),
       .io_b_4( io_y_4 ),
       .io_b_3( io_y_3 ),
       .io_b_2( io_y_2 ),
       .io_b_1( io_y_1 ),
       .io_b_0( io_y_0 ),
       .io_o_2( MatrixVectorMultModule_io_o_2 ),
       .io_o_1( MatrixVectorMultModule_io_o_1 ),
       .io_o_0( MatrixVectorMultModule_io_o_0 )
  );
  MatrixVectorMultModule_0 MatrixVectorMultModule_1(.clk(clk),
       .io_a_2_2( io_c_2_2 ),
       .io_a_2_1( io_c_1_2 ),
       .io_a_2_0( io_c_0_2 ),
       .io_a_1_2( io_c_2_1 ),
       .io_a_1_1( io_c_1_1 ),
       .io_a_1_0( io_c_0_1 ),
       .io_a_0_2( io_c_2_0 ),
       .io_a_0_1( io_c_1_0 ),
       .io_a_0_0( io_c_0_0 ),
       .io_b_2( io_z_2 ),
       .io_b_1( io_z_1 ),
       .io_b_0( io_z_0 ),
       .io_o_2( MatrixVectorMultModule_1_io_o_2 ),
       .io_o_1( MatrixVectorMultModule_1_io_o_1 ),
       .io_o_0( MatrixVectorMultModule_1_io_o_0 )
  );
  gModule gModule(
       .io_in( x_stage_0 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_io_ou )
  );
  gModule gModule_1(
       .io_in( x_stage_1 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_1_io_ou )
  );
  gModule gModule_2(
       .io_in( x_stage_2 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_2_io_ou )
  );

  always @(posedge clk) begin
    x_stage_2 <= T0;
    cz_2 <= MatrixVectorMultModule_1_io_o_2;
    xay_2 <= T4;
    x_delay_2 <= R8;
    R8 <= io_x_2;
    x_stage_1 <= T9;
    cz_1 <= MatrixVectorMultModule_1_io_o_1;
    xay_1 <= T13;
    x_delay_1 <= R17;
    R17 <= io_x_1;
    x_stage_0 <= T18;
    cz_0 <= MatrixVectorMultModule_1_io_o_0;
    xay_0 <= T22;
    x_delay_0 <= R26;
    R26 <= io_x_0;
  end
endmodule

module MatrixVectorMultModule_2(input clk,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    output[17:0] io_o_11,
    output[17:0] io_o_10,
    output[17:0] io_o_9,
    output[17:0] io_o_8,
    output[17:0] io_o_7,
    output[17:0] io_o_6,
    output[17:0] io_o_5,
    output[17:0] io_o_4,
    output[17:0] io_o_3,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] R0;
  reg [17:0] R1;
  reg [17:0] R2;
  reg [17:0] R3;
  reg [17:0] R4;
  reg [17:0] R5;
  reg [17:0] R6;
  reg [17:0] R7;
  reg [17:0] R8;
  reg [17:0] R9;
  reg [17:0] R10;
  reg [17:0] R11;
  wire[17:0] DotProductModule_io_o;
  wire[17:0] DotProductModule_1_io_o;
  wire[17:0] DotProductModule_2_io_o;
  wire[17:0] DotProductModule_3_io_o;
  wire[17:0] DotProductModule_4_io_o;
  wire[17:0] DotProductModule_5_io_o;
  wire[17:0] DotProductModule_6_io_o;
  wire[17:0] DotProductModule_7_io_o;
  wire[17:0] DotProductModule_8_io_o;
  wire[17:0] DotProductModule_9_io_o;
  wire[17:0] DotProductModule_10_io_o;
  wire[17:0] DotProductModule_11_io_o;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
    R2 = {1{$random}};
    R3 = {1{$random}};
    R4 = {1{$random}};
    R5 = {1{$random}};
    R6 = {1{$random}};
    R7 = {1{$random}};
    R8 = {1{$random}};
    R9 = {1{$random}};
    R10 = {1{$random}};
    R11 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_o_0 = R0;
  assign io_o_1 = R1;
  assign io_o_2 = R2;
  assign io_o_3 = R3;
  assign io_o_4 = R4;
  assign io_o_5 = R5;
  assign io_o_6 = R6;
  assign io_o_7 = R7;
  assign io_o_8 = R8;
  assign io_o_9 = R9;
  assign io_o_10 = R10;
  assign io_o_11 = R11;
  DotProductModule_0 DotProductModule(.clk(clk),
       .io_a_2( io_a_0_2 ),
       .io_a_1( io_a_0_1 ),
       .io_a_0( io_a_0_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_io_o )
  );
  DotProductModule_0 DotProductModule_1(.clk(clk),
       .io_a_2( io_a_1_2 ),
       .io_a_1( io_a_1_1 ),
       .io_a_0( io_a_1_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_1_io_o )
  );
  DotProductModule_0 DotProductModule_2(.clk(clk),
       .io_a_2( io_a_2_2 ),
       .io_a_1( io_a_2_1 ),
       .io_a_0( io_a_2_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_2_io_o )
  );
  DotProductModule_0 DotProductModule_3(.clk(clk),
       .io_a_2( io_a_3_2 ),
       .io_a_1( io_a_3_1 ),
       .io_a_0( io_a_3_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_3_io_o )
  );
  DotProductModule_0 DotProductModule_4(.clk(clk),
       .io_a_2( io_a_4_2 ),
       .io_a_1( io_a_4_1 ),
       .io_a_0( io_a_4_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_4_io_o )
  );
  DotProductModule_0 DotProductModule_5(.clk(clk),
       .io_a_2( io_a_5_2 ),
       .io_a_1( io_a_5_1 ),
       .io_a_0( io_a_5_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_5_io_o )
  );
  DotProductModule_0 DotProductModule_6(.clk(clk),
       .io_a_2( io_a_6_2 ),
       .io_a_1( io_a_6_1 ),
       .io_a_0( io_a_6_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_6_io_o )
  );
  DotProductModule_0 DotProductModule_7(.clk(clk),
       .io_a_2( io_a_7_2 ),
       .io_a_1( io_a_7_1 ),
       .io_a_0( io_a_7_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_7_io_o )
  );
  DotProductModule_0 DotProductModule_8(.clk(clk),
       .io_a_2( io_a_8_2 ),
       .io_a_1( io_a_8_1 ),
       .io_a_0( io_a_8_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_8_io_o )
  );
  DotProductModule_0 DotProductModule_9(.clk(clk),
       .io_a_2( io_a_9_2 ),
       .io_a_1( io_a_9_1 ),
       .io_a_0( io_a_9_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_9_io_o )
  );
  DotProductModule_0 DotProductModule_10(.clk(clk),
       .io_a_2( io_a_10_2 ),
       .io_a_1( io_a_10_1 ),
       .io_a_0( io_a_10_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_10_io_o )
  );
  DotProductModule_0 DotProductModule_11(.clk(clk),
       .io_a_2( io_a_11_2 ),
       .io_a_1( io_a_11_1 ),
       .io_a_0( io_a_11_0 ),
       .io_b_2( io_b_2 ),
       .io_b_1( io_b_1 ),
       .io_b_0( io_b_0 ),
       .io_o( DotProductModule_11_io_o )
  );

  always @(posedge clk) begin
    R0 <= DotProductModule_io_o;
    R1 <= DotProductModule_1_io_o;
    R2 <= DotProductModule_2_io_o;
    R3 <= DotProductModule_3_io_o;
    R4 <= DotProductModule_4_io_o;
    R5 <= DotProductModule_5_io_o;
    R6 <= DotProductModule_6_io_o;
    R7 <= DotProductModule_7_io_o;
    R8 <= DotProductModule_8_io_o;
    R9 <= DotProductModule_9_io_o;
    R10 <= DotProductModule_10_io_o;
    R11 <= DotProductModule_11_io_o;
  end
endmodule

module YNetModule(input clk,
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_y_11,
    input [17:0] io_y_10,
    input [17:0] io_y_9,
    input [17:0] io_y_8,
    input [17:0] io_y_7,
    input [17:0] io_y_6,
    input [17:0] io_y_5,
    input [17:0] io_y_4,
    input [17:0] io_y_3,
    input [17:0] io_y_2,
    input [17:0] io_y_1,
    input [17:0] io_y_0,
    input [17:0] io_b_11,
    input [17:0] io_b_10,
    input [17:0] io_b_9,
    input [17:0] io_b_8,
    input [17:0] io_b_7,
    input [17:0] io_b_6,
    input [17:0] io_b_5,
    input [17:0] io_b_4,
    input [17:0] io_b_3,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    output[17:0] io_o_11,
    output[17:0] io_o_10,
    output[17:0] io_o_9,
    output[17:0] io_o_8,
    output[17:0] io_o_7,
    output[17:0] io_o_6,
    output[17:0] io_o_5,
    output[17:0] io_o_4,
    output[17:0] io_o_3,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] y_stage_11;
  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  reg [17:0] y_next_11;
  reg [17:0] R3;
  reg [17:0] R4;
  wire[17:0] T5;
  reg [17:0] axb_11;
  wire[17:0] T6;
  wire[17:0] T7;
  wire[17:0] T8;
  reg [17:0] b_next_11;
  reg [17:0] R9;
  wire[17:0] T10;
  reg [17:0] y_stage_10;
  wire[17:0] T11;
  wire[17:0] T12;
  wire[17:0] T13;
  reg [17:0] y_next_10;
  reg [17:0] R14;
  reg [17:0] R15;
  wire[17:0] T16;
  reg [17:0] axb_10;
  wire[17:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  reg [17:0] b_next_10;
  reg [17:0] R20;
  wire[17:0] T21;
  reg [17:0] y_stage_9;
  wire[17:0] T22;
  wire[17:0] T23;
  wire[17:0] T24;
  reg [17:0] y_next_9;
  reg [17:0] R25;
  reg [17:0] R26;
  wire[17:0] T27;
  reg [17:0] axb_9;
  wire[17:0] T28;
  wire[17:0] T29;
  wire[17:0] T30;
  reg [17:0] b_next_9;
  reg [17:0] R31;
  wire[17:0] T32;
  reg [17:0] y_stage_8;
  wire[17:0] T33;
  wire[17:0] T34;
  wire[17:0] T35;
  reg [17:0] y_next_8;
  reg [17:0] R36;
  reg [17:0] R37;
  wire[17:0] T38;
  reg [17:0] axb_8;
  wire[17:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  reg [17:0] b_next_8;
  reg [17:0] R42;
  wire[17:0] T43;
  reg [17:0] y_stage_7;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[17:0] T46;
  reg [17:0] y_next_7;
  reg [17:0] R47;
  reg [17:0] R48;
  wire[17:0] T49;
  reg [17:0] axb_7;
  wire[17:0] T50;
  wire[17:0] T51;
  wire[17:0] T52;
  reg [17:0] b_next_7;
  reg [17:0] R53;
  wire[17:0] T54;
  reg [17:0] y_stage_6;
  wire[17:0] T55;
  wire[17:0] T56;
  wire[17:0] T57;
  reg [17:0] y_next_6;
  reg [17:0] R58;
  reg [17:0] R59;
  wire[17:0] T60;
  reg [17:0] axb_6;
  wire[17:0] T61;
  wire[17:0] T62;
  wire[17:0] T63;
  reg [17:0] b_next_6;
  reg [17:0] R64;
  wire[17:0] T65;
  reg [17:0] y_stage_5;
  wire[17:0] T66;
  wire[17:0] T67;
  wire[17:0] T68;
  reg [17:0] y_next_5;
  reg [17:0] R69;
  reg [17:0] R70;
  wire[17:0] T71;
  reg [17:0] axb_5;
  wire[17:0] T72;
  wire[17:0] T73;
  wire[17:0] T74;
  reg [17:0] b_next_5;
  reg [17:0] R75;
  wire[17:0] T76;
  reg [17:0] y_stage_4;
  wire[17:0] T77;
  wire[17:0] T78;
  wire[17:0] T79;
  reg [17:0] y_next_4;
  reg [17:0] R80;
  reg [17:0] R81;
  wire[17:0] T82;
  reg [17:0] axb_4;
  wire[17:0] T83;
  wire[17:0] T84;
  wire[17:0] T85;
  reg [17:0] b_next_4;
  reg [17:0] R86;
  wire[17:0] T87;
  reg [17:0] y_stage_3;
  wire[17:0] T88;
  wire[17:0] T89;
  wire[17:0] T90;
  reg [17:0] y_next_3;
  reg [17:0] R91;
  reg [17:0] R92;
  wire[17:0] T93;
  reg [17:0] axb_3;
  wire[17:0] T94;
  wire[17:0] T95;
  wire[17:0] T96;
  reg [17:0] b_next_3;
  reg [17:0] R97;
  wire[17:0] T98;
  reg [17:0] y_stage_2;
  wire[17:0] T99;
  wire[17:0] T100;
  wire[17:0] T101;
  reg [17:0] y_next_2;
  reg [17:0] R102;
  reg [17:0] R103;
  wire[17:0] T104;
  reg [17:0] axb_2;
  wire[17:0] T105;
  wire[17:0] T106;
  wire[17:0] T107;
  reg [17:0] b_next_2;
  reg [17:0] R108;
  wire[17:0] T109;
  reg [17:0] y_stage_1;
  wire[17:0] T110;
  wire[17:0] T111;
  wire[17:0] T112;
  reg [17:0] y_next_1;
  reg [17:0] R113;
  reg [17:0] R114;
  wire[17:0] T115;
  reg [17:0] axb_1;
  wire[17:0] T116;
  wire[17:0] T117;
  wire[17:0] T118;
  reg [17:0] b_next_1;
  reg [17:0] R119;
  wire[17:0] T120;
  reg [17:0] y_stage_0;
  wire[17:0] T121;
  wire[17:0] T122;
  wire[17:0] T123;
  reg [17:0] y_next_0;
  reg [17:0] R124;
  reg [17:0] R125;
  wire[17:0] T126;
  reg [17:0] axb_0;
  wire[17:0] T127;
  wire[17:0] T128;
  wire[17:0] T129;
  reg [17:0] b_next_0;
  reg [17:0] R130;
  wire[17:0] T131;
  wire[17:0] gModule_io_ou;
  wire[17:0] gModule_1_io_ou;
  wire[17:0] gModule_2_io_ou;
  wire[17:0] gModule_3_io_ou;
  wire[17:0] gModule_4_io_ou;
  wire[17:0] gModule_5_io_ou;
  wire[17:0] gModule_6_io_ou;
  wire[17:0] gModule_7_io_ou;
  wire[17:0] gModule_8_io_ou;
  wire[17:0] gModule_9_io_ou;
  wire[17:0] gModule_10_io_ou;
  wire[17:0] gModule_11_io_ou;
  wire[17:0] MatrixVectorMultModule_io_o_11;
  wire[17:0] MatrixVectorMultModule_io_o_10;
  wire[17:0] MatrixVectorMultModule_io_o_9;
  wire[17:0] MatrixVectorMultModule_io_o_8;
  wire[17:0] MatrixVectorMultModule_io_o_7;
  wire[17:0] MatrixVectorMultModule_io_o_6;
  wire[17:0] MatrixVectorMultModule_io_o_5;
  wire[17:0] MatrixVectorMultModule_io_o_4;
  wire[17:0] MatrixVectorMultModule_io_o_3;
  wire[17:0] MatrixVectorMultModule_io_o_2;
  wire[17:0] MatrixVectorMultModule_io_o_1;
  wire[17:0] MatrixVectorMultModule_io_o_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    y_stage_11 = {1{$random}};
    y_next_11 = {1{$random}};
    R3 = {1{$random}};
    R4 = {1{$random}};
    axb_11 = {1{$random}};
    b_next_11 = {1{$random}};
    R9 = {1{$random}};
    y_stage_10 = {1{$random}};
    y_next_10 = {1{$random}};
    R14 = {1{$random}};
    R15 = {1{$random}};
    axb_10 = {1{$random}};
    b_next_10 = {1{$random}};
    R20 = {1{$random}};
    y_stage_9 = {1{$random}};
    y_next_9 = {1{$random}};
    R25 = {1{$random}};
    R26 = {1{$random}};
    axb_9 = {1{$random}};
    b_next_9 = {1{$random}};
    R31 = {1{$random}};
    y_stage_8 = {1{$random}};
    y_next_8 = {1{$random}};
    R36 = {1{$random}};
    R37 = {1{$random}};
    axb_8 = {1{$random}};
    b_next_8 = {1{$random}};
    R42 = {1{$random}};
    y_stage_7 = {1{$random}};
    y_next_7 = {1{$random}};
    R47 = {1{$random}};
    R48 = {1{$random}};
    axb_7 = {1{$random}};
    b_next_7 = {1{$random}};
    R53 = {1{$random}};
    y_stage_6 = {1{$random}};
    y_next_6 = {1{$random}};
    R58 = {1{$random}};
    R59 = {1{$random}};
    axb_6 = {1{$random}};
    b_next_6 = {1{$random}};
    R64 = {1{$random}};
    y_stage_5 = {1{$random}};
    y_next_5 = {1{$random}};
    R69 = {1{$random}};
    R70 = {1{$random}};
    axb_5 = {1{$random}};
    b_next_5 = {1{$random}};
    R75 = {1{$random}};
    y_stage_4 = {1{$random}};
    y_next_4 = {1{$random}};
    R80 = {1{$random}};
    R81 = {1{$random}};
    axb_4 = {1{$random}};
    b_next_4 = {1{$random}};
    R86 = {1{$random}};
    y_stage_3 = {1{$random}};
    y_next_3 = {1{$random}};
    R91 = {1{$random}};
    R92 = {1{$random}};
    axb_3 = {1{$random}};
    b_next_3 = {1{$random}};
    R97 = {1{$random}};
    y_stage_2 = {1{$random}};
    y_next_2 = {1{$random}};
    R102 = {1{$random}};
    R103 = {1{$random}};
    axb_2 = {1{$random}};
    b_next_2 = {1{$random}};
    R108 = {1{$random}};
    y_stage_1 = {1{$random}};
    y_next_1 = {1{$random}};
    R113 = {1{$random}};
    R114 = {1{$random}};
    axb_1 = {1{$random}};
    b_next_1 = {1{$random}};
    R119 = {1{$random}};
    y_stage_0 = {1{$random}};
    y_next_0 = {1{$random}};
    R124 = {1{$random}};
    R125 = {1{$random}};
    axb_0 = {1{$random}};
    b_next_0 = {1{$random}};
    R130 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T1;
  assign T1 = T5 + T2;
  assign T2 = y_next_11;
  assign T5 = axb_11;
  assign T6 = T7;
  assign T7 = T10 - T8;
  assign T8 = b_next_11;
  assign T10 = MatrixVectorMultModule_io_o_11;
  assign T11 = T12;
  assign T12 = T16 + T13;
  assign T13 = y_next_10;
  assign T16 = axb_10;
  assign T17 = T18;
  assign T18 = T21 - T19;
  assign T19 = b_next_10;
  assign T21 = MatrixVectorMultModule_io_o_10;
  assign T22 = T23;
  assign T23 = T27 + T24;
  assign T24 = y_next_9;
  assign T27 = axb_9;
  assign T28 = T29;
  assign T29 = T32 - T30;
  assign T30 = b_next_9;
  assign T32 = MatrixVectorMultModule_io_o_9;
  assign T33 = T34;
  assign T34 = T38 + T35;
  assign T35 = y_next_8;
  assign T38 = axb_8;
  assign T39 = T40;
  assign T40 = T43 - T41;
  assign T41 = b_next_8;
  assign T43 = MatrixVectorMultModule_io_o_8;
  assign T44 = T45;
  assign T45 = T49 + T46;
  assign T46 = y_next_7;
  assign T49 = axb_7;
  assign T50 = T51;
  assign T51 = T54 - T52;
  assign T52 = b_next_7;
  assign T54 = MatrixVectorMultModule_io_o_7;
  assign T55 = T56;
  assign T56 = T60 + T57;
  assign T57 = y_next_6;
  assign T60 = axb_6;
  assign T61 = T62;
  assign T62 = T65 - T63;
  assign T63 = b_next_6;
  assign T65 = MatrixVectorMultModule_io_o_6;
  assign T66 = T67;
  assign T67 = T71 + T68;
  assign T68 = y_next_5;
  assign T71 = axb_5;
  assign T72 = T73;
  assign T73 = T76 - T74;
  assign T74 = b_next_5;
  assign T76 = MatrixVectorMultModule_io_o_5;
  assign T77 = T78;
  assign T78 = T82 + T79;
  assign T79 = y_next_4;
  assign T82 = axb_4;
  assign T83 = T84;
  assign T84 = T87 - T85;
  assign T85 = b_next_4;
  assign T87 = MatrixVectorMultModule_io_o_4;
  assign T88 = T89;
  assign T89 = T93 + T90;
  assign T90 = y_next_3;
  assign T93 = axb_3;
  assign T94 = T95;
  assign T95 = T98 - T96;
  assign T96 = b_next_3;
  assign T98 = MatrixVectorMultModule_io_o_3;
  assign T99 = T100;
  assign T100 = T104 + T101;
  assign T101 = y_next_2;
  assign T104 = axb_2;
  assign T105 = T106;
  assign T106 = T109 - T107;
  assign T107 = b_next_2;
  assign T109 = MatrixVectorMultModule_io_o_2;
  assign T110 = T111;
  assign T111 = T115 + T112;
  assign T112 = y_next_1;
  assign T115 = axb_1;
  assign T116 = T117;
  assign T117 = T120 - T118;
  assign T118 = b_next_1;
  assign T120 = MatrixVectorMultModule_io_o_1;
  assign T121 = T122;
  assign T122 = T126 + T123;
  assign T123 = y_next_0;
  assign T126 = axb_0;
  assign T127 = T128;
  assign T128 = T131 - T129;
  assign T129 = b_next_0;
  assign T131 = MatrixVectorMultModule_io_o_0;
  assign io_o_0 = gModule_io_ou;
  assign io_o_1 = gModule_1_io_ou;
  assign io_o_2 = gModule_2_io_ou;
  assign io_o_3 = gModule_3_io_ou;
  assign io_o_4 = gModule_4_io_ou;
  assign io_o_5 = gModule_5_io_ou;
  assign io_o_6 = gModule_6_io_ou;
  assign io_o_7 = gModule_7_io_ou;
  assign io_o_8 = gModule_8_io_ou;
  assign io_o_9 = gModule_9_io_ou;
  assign io_o_10 = gModule_10_io_ou;
  assign io_o_11 = gModule_11_io_ou;
  MatrixVectorMultModule_2 MatrixVectorMultModule(.clk(clk),
       .io_a_11_2( io_a_11_2 ),
       .io_a_11_1( io_a_11_1 ),
       .io_a_11_0( io_a_11_0 ),
       .io_a_10_2( io_a_10_2 ),
       .io_a_10_1( io_a_10_1 ),
       .io_a_10_0( io_a_10_0 ),
       .io_a_9_2( io_a_9_2 ),
       .io_a_9_1( io_a_9_1 ),
       .io_a_9_0( io_a_9_0 ),
       .io_a_8_2( io_a_8_2 ),
       .io_a_8_1( io_a_8_1 ),
       .io_a_8_0( io_a_8_0 ),
       .io_a_7_2( io_a_7_2 ),
       .io_a_7_1( io_a_7_1 ),
       .io_a_7_0( io_a_7_0 ),
       .io_a_6_2( io_a_6_2 ),
       .io_a_6_1( io_a_6_1 ),
       .io_a_6_0( io_a_6_0 ),
       .io_a_5_2( io_a_5_2 ),
       .io_a_5_1( io_a_5_1 ),
       .io_a_5_0( io_a_5_0 ),
       .io_a_4_2( io_a_4_2 ),
       .io_a_4_1( io_a_4_1 ),
       .io_a_4_0( io_a_4_0 ),
       .io_a_3_2( io_a_3_2 ),
       .io_a_3_1( io_a_3_1 ),
       .io_a_3_0( io_a_3_0 ),
       .io_a_2_2( io_a_2_2 ),
       .io_a_2_1( io_a_2_1 ),
       .io_a_2_0( io_a_2_0 ),
       .io_a_1_2( io_a_1_2 ),
       .io_a_1_1( io_a_1_1 ),
       .io_a_1_0( io_a_1_0 ),
       .io_a_0_2( io_a_0_2 ),
       .io_a_0_1( io_a_0_1 ),
       .io_a_0_0( io_a_0_0 ),
       .io_b_2( io_x_2 ),
       .io_b_1( io_x_1 ),
       .io_b_0( io_x_0 ),
       .io_o_11( MatrixVectorMultModule_io_o_11 ),
       .io_o_10( MatrixVectorMultModule_io_o_10 ),
       .io_o_9( MatrixVectorMultModule_io_o_9 ),
       .io_o_8( MatrixVectorMultModule_io_o_8 ),
       .io_o_7( MatrixVectorMultModule_io_o_7 ),
       .io_o_6( MatrixVectorMultModule_io_o_6 ),
       .io_o_5( MatrixVectorMultModule_io_o_5 ),
       .io_o_4( MatrixVectorMultModule_io_o_4 ),
       .io_o_3( MatrixVectorMultModule_io_o_3 ),
       .io_o_2( MatrixVectorMultModule_io_o_2 ),
       .io_o_1( MatrixVectorMultModule_io_o_1 ),
       .io_o_0( MatrixVectorMultModule_io_o_0 )
  );
  gModule gModule(
       .io_in( y_stage_0 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_io_ou )
  );
  gModule gModule_1(
       .io_in( y_stage_1 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_1_io_ou )
  );
  gModule gModule_2(
       .io_in( y_stage_2 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_2_io_ou )
  );
  gModule gModule_3(
       .io_in( y_stage_3 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_3_io_ou )
  );
  gModule gModule_4(
       .io_in( y_stage_4 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_4_io_ou )
  );
  gModule gModule_5(
       .io_in( y_stage_5 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_5_io_ou )
  );
  gModule gModule_6(
       .io_in( y_stage_6 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_6_io_ou )
  );
  gModule gModule_7(
       .io_in( y_stage_7 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_7_io_ou )
  );
  gModule gModule_8(
       .io_in( y_stage_8 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_8_io_ou )
  );
  gModule gModule_9(
       .io_in( y_stage_9 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_9_io_ou )
  );
  gModule gModule_10(
       .io_in( y_stage_10 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_10_io_ou )
  );
  gModule gModule_11(
       .io_in( y_stage_11 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_11_io_ou )
  );

  always @(posedge clk) begin
    y_stage_11 <= T0;
    y_next_11 <= R3;
    R3 <= R4;
    R4 <= io_y_11;
    axb_11 <= T6;
    b_next_11 <= R9;
    R9 <= io_b_11;
    y_stage_10 <= T11;
    y_next_10 <= R14;
    R14 <= R15;
    R15 <= io_y_10;
    axb_10 <= T17;
    b_next_10 <= R20;
    R20 <= io_b_10;
    y_stage_9 <= T22;
    y_next_9 <= R25;
    R25 <= R26;
    R26 <= io_y_9;
    axb_9 <= T28;
    b_next_9 <= R31;
    R31 <= io_b_9;
    y_stage_8 <= T33;
    y_next_8 <= R36;
    R36 <= R37;
    R37 <= io_y_8;
    axb_8 <= T39;
    b_next_8 <= R42;
    R42 <= io_b_8;
    y_stage_7 <= T44;
    y_next_7 <= R47;
    R47 <= R48;
    R48 <= io_y_7;
    axb_7 <= T50;
    b_next_7 <= R53;
    R53 <= io_b_7;
    y_stage_6 <= T55;
    y_next_6 <= R58;
    R58 <= R59;
    R59 <= io_y_6;
    axb_6 <= T61;
    b_next_6 <= R64;
    R64 <= io_b_6;
    y_stage_5 <= T66;
    y_next_5 <= R69;
    R69 <= R70;
    R70 <= io_y_5;
    axb_5 <= T72;
    b_next_5 <= R75;
    R75 <= io_b_5;
    y_stage_4 <= T77;
    y_next_4 <= R80;
    R80 <= R81;
    R81 <= io_y_4;
    axb_4 <= T83;
    b_next_4 <= R86;
    R86 <= io_b_4;
    y_stage_3 <= T88;
    y_next_3 <= R91;
    R91 <= R92;
    R92 <= io_y_3;
    axb_3 <= T94;
    b_next_3 <= R97;
    R97 <= io_b_3;
    y_stage_2 <= T99;
    y_next_2 <= R102;
    R102 <= R103;
    R103 <= io_y_2;
    axb_2 <= T105;
    b_next_2 <= R108;
    R108 <= io_b_2;
    y_stage_1 <= T110;
    y_next_1 <= R113;
    R113 <= R114;
    R114 <= io_y_1;
    axb_1 <= T116;
    b_next_1 <= R119;
    R119 <= io_b_1;
    y_stage_0 <= T121;
    y_next_0 <= R124;
    R124 <= R125;
    R125 <= io_y_0;
    axb_0 <= T127;
    b_next_0 <= R130;
    R130 <= io_b_0;
  end
endmodule

module ZNetModule(input clk,
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_z_2,
    input [17:0] io_z_1,
    input [17:0] io_z_0,
    input [17:0] io_c_2_2,
    input [17:0] io_c_2_1,
    input [17:0] io_c_2_0,
    input [17:0] io_c_1_2,
    input [17:0] io_c_1_1,
    input [17:0] io_c_1_0,
    input [17:0] io_c_0_2,
    input [17:0] io_c_0_1,
    input [17:0] io_c_0_0,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  reg [17:0] z_stage_2;
  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  reg [17:0] z_next_2;
  reg [17:0] R3;
  wire[17:0] T4;
  reg [17:0] z_stage_1;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  reg [17:0] z_next_1;
  reg [17:0] R8;
  wire[17:0] T9;
  reg [17:0] z_stage_0;
  wire[17:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  reg [17:0] z_next_0;
  reg [17:0] R13;
  wire[17:0] T14;
  wire[17:0] gModule_io_ou;
  wire[17:0] gModule_1_io_ou;
  wire[17:0] gModule_2_io_ou;
  wire[17:0] MatrixVectorMultModule_io_o_2;
  wire[17:0] MatrixVectorMultModule_io_o_1;
  wire[17:0] MatrixVectorMultModule_io_o_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    z_stage_2 = {1{$random}};
    z_next_2 = {1{$random}};
    R3 = {1{$random}};
    z_stage_1 = {1{$random}};
    z_next_1 = {1{$random}};
    R8 = {1{$random}};
    z_stage_0 = {1{$random}};
    z_next_0 = {1{$random}};
    R13 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T1;
  assign T1 = T4 - T2;
  assign T2 = z_next_2;
  assign T4 = MatrixVectorMultModule_io_o_2;
  assign T5 = T6;
  assign T6 = T9 - T7;
  assign T7 = z_next_1;
  assign T9 = MatrixVectorMultModule_io_o_1;
  assign T10 = T11;
  assign T11 = T14 - T12;
  assign T12 = z_next_0;
  assign T14 = MatrixVectorMultModule_io_o_0;
  assign io_o_0 = gModule_io_ou;
  assign io_o_1 = gModule_1_io_ou;
  assign io_o_2 = gModule_2_io_ou;
  MatrixVectorMultModule_0 MatrixVectorMultModule(.clk(clk),
       .io_a_2_2( io_c_2_2 ),
       .io_a_2_1( io_c_2_1 ),
       .io_a_2_0( io_c_2_0 ),
       .io_a_1_2( io_c_1_2 ),
       .io_a_1_1( io_c_1_1 ),
       .io_a_1_0( io_c_1_0 ),
       .io_a_0_2( io_c_0_2 ),
       .io_a_0_1( io_c_0_1 ),
       .io_a_0_0( io_c_0_0 ),
       .io_b_2( io_x_2 ),
       .io_b_1( io_x_1 ),
       .io_b_0( io_x_0 ),
       .io_o_2( MatrixVectorMultModule_io_o_2 ),
       .io_o_1( MatrixVectorMultModule_io_o_1 ),
       .io_o_0( MatrixVectorMultModule_io_o_0 )
  );
  gModule gModule(
       .io_in( z_stage_0 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_io_ou )
  );
  gModule gModule_1(
       .io_in( z_stage_1 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_1_io_ou )
  );
  gModule gModule_2(
       .io_in( z_stage_2 ),
       .io_hi( 18'h8000 ),
       .io_lo( 18'h38000 ),
       .io_ou( gModule_2_io_ou )
  );

  always @(posedge clk) begin
    z_stage_2 <= T0;
    z_next_2 <= R3;
    R3 <= io_z_2;
    z_stage_1 <= T5;
    z_next_1 <= R8;
    R8 <= io_z_1;
    z_stage_0 <= T10;
    z_next_0 <= R13;
    R13 <= io_z_0;
  end
endmodule

module NN1Top(input clk,
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_y_11,
    input [17:0] io_y_10,
    input [17:0] io_y_9,
    input [17:0] io_y_8,
    input [17:0] io_y_7,
    input [17:0] io_y_6,
    input [17:0] io_y_5,
    input [17:0] io_y_4,
    input [17:0] io_y_3,
    input [17:0] io_y_2,
    input [17:0] io_y_1,
    input [17:0] io_y_0,
    input [17:0] io_z_2,
    input [17:0] io_z_1,
    input [17:0] io_z_0,
    input [17:0] io_b_11,
    input [17:0] io_b_10,
    input [17:0] io_b_9,
    input [17:0] io_b_8,
    input [17:0] io_b_7,
    input [17:0] io_b_6,
    input [17:0] io_b_5,
    input [17:0] io_b_4,
    input [17:0] io_b_3,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_c_2_2,
    input [17:0] io_c_2_1,
    input [17:0] io_c_2_0,
    input [17:0] io_c_1_2,
    input [17:0] io_c_1_1,
    input [17:0] io_c_1_0,
    input [17:0] io_c_0_2,
    input [17:0] io_c_0_1,
    input [17:0] io_c_0_0,
    input [17:0] io_lbda,
    output[17:0] io_xout_2,
    output[17:0] io_xout_1,
    output[17:0] io_xout_0,
    output[17:0] io_yout_11,
    output[17:0] io_yout_10,
    output[17:0] io_yout_9,
    output[17:0] io_yout_8,
    output[17:0] io_yout_7,
    output[17:0] io_yout_6,
    output[17:0] io_yout_5,
    output[17:0] io_yout_4,
    output[17:0] io_yout_3,
    output[17:0] io_yout_2,
    output[17:0] io_yout_1,
    output[17:0] io_yout_0,
    output[17:0] io_zout_2,
    output[17:0] io_zout_1,
    output[17:0] io_zout_0
);

  reg [17:0] R0;
  reg [17:0] R1;
  reg [17:0] R2;
  reg [17:0] R3;
  reg [17:0] R4;
  reg [17:0] R5;
  reg [17:0] R6;
  reg [17:0] R7;
  reg [17:0] R8;
  reg [17:0] R9;
  reg [17:0] R10;
  reg [17:0] R11;
  reg [17:0] R12;
  reg [17:0] R13;
  reg [17:0] R14;
  reg [17:0] R15;
  reg [17:0] R16;
  reg [17:0] R17;
  reg [17:0] R18;
  reg [17:0] R19;
  reg [17:0] R20;
  reg [17:0] R21;
  reg [17:0] R22;
  reg [17:0] R23;
  reg [17:0] R24;
  reg [17:0] R25;
  reg [17:0] R26;
  reg [17:0] R27;
  reg [17:0] R28;
  reg [17:0] R29;
  reg [17:0] R30;
  reg [17:0] R31;
  reg [17:0] R32;
  reg [17:0] R33;
  reg [17:0] R34;
  reg [17:0] R35;
  reg [17:0] R36;
  reg [17:0] R37;
  reg [17:0] R38;
  reg [17:0] R39;
  reg [17:0] R40;
  reg [17:0] R41;
  reg [17:0] R42;
  reg [17:0] R43;
  reg [17:0] R44;
  reg [17:0] R45;
  reg [17:0] R46;
  reg [17:0] R47;
  reg [17:0] R48;
  reg [17:0] R49;
  reg [17:0] R50;
  reg [17:0] R51;
  reg [17:0] R52;
  reg [17:0] R53;
  reg [17:0] R54;
  reg [17:0] R55;
  reg [17:0] R56;
  reg [17:0] R57;
  reg [17:0] R58;
  reg [17:0] R59;
  reg [17:0] R60;
  reg [17:0] R61;
  reg [17:0] R62;
  reg [17:0] R63;
  reg [17:0] R64;
  reg [17:0] R65;
  reg [17:0] R66;
  reg [17:0] R67;
  reg [17:0] R68;
  reg [17:0] R69;
  reg [17:0] R70;
  reg [17:0] R71;
  reg [17:0] R72;
  reg [17:0] R73;
  reg [17:0] R74;
  reg [17:0] R75;
  reg [17:0] R76;
  reg [17:0] R77;
  reg [17:0] R78;
  reg [17:0] R79;
  reg [17:0] R80;
  reg [17:0] R81;
  reg [17:0] R82;
  reg [17:0] R83;
  reg [17:0] R84;
  reg [17:0] R85;
  reg [17:0] R86;
  reg [17:0] R87;
  reg [17:0] R88;
  reg [17:0] R89;
  reg [17:0] R90;
  reg [17:0] R91;
  reg [17:0] R92;
  reg [17:0] R93;
  reg [17:0] R94;
  reg [17:0] R95;
  reg [17:0] R96;
  reg [17:0] R97;
  reg [17:0] R98;
  reg [17:0] R99;
  reg [17:0] R100;
  reg [17:0] R101;
  reg [17:0] R102;
  reg [17:0] R103;
  reg [17:0] R104;
  reg [17:0] R105;
  reg [17:0] R106;
  reg [17:0] R107;
  reg [17:0] R108;
  reg [17:0] R109;
  reg [17:0] R110;
  reg [17:0] R111;
  reg [17:0] R112;
  reg [17:0] R113;
  reg [17:0] R114;
  reg [17:0] R115;
  reg [17:0] R116;
  reg [17:0] R117;
  reg [17:0] R118;
  reg [17:0] R119;
  reg [17:0] R120;
  reg [17:0] R121;
  reg [17:0] R122;
  reg [17:0] R123;
  reg [17:0] R124;
  reg [17:0] R125;
  reg [17:0] R126;
  reg [17:0] R127;
  reg [17:0] R128;
  reg [17:0] R129;
  reg [17:0] R130;
  reg [17:0] R131;
  reg [17:0] R132;
  reg [17:0] R133;
  reg [17:0] R134;
  reg [17:0] R135;
  reg [17:0] R136;
  reg [17:0] R137;
  reg [17:0] R138;
  reg [17:0] R139;
  reg [17:0] R140;
  reg [17:0] R141;
  reg [17:0] R142;
  reg [17:0] R143;
  reg [17:0] R144;
  reg [17:0] R145;
  reg [17:0] R146;
  reg [17:0] R147;
  reg [17:0] R148;
  reg [17:0] R149;
  reg [17:0] R150;
  reg [17:0] R151;
  reg [17:0] R152;
  reg [17:0] R153;
  reg [17:0] R154;
  reg [17:0] R155;
  reg [17:0] R156;
  reg [17:0] R157;
  reg [17:0] R158;
  reg [17:0] R159;
  reg [17:0] R160;
  reg [17:0] R161;
  reg [17:0] R162;
  reg [17:0] R163;
  reg [17:0] R164;
  reg [17:0] R165;
  reg [17:0] R166;
  reg [17:0] R167;
  reg [17:0] R168;
  reg [17:0] R169;
  reg [17:0] R170;
  reg [17:0] R171;
  reg [17:0] R172;
  reg [17:0] R173;
  reg [17:0] R174;
  reg [17:0] R175;
  reg [17:0] R176;
  reg [17:0] R177;
  reg [17:0] R178;
  reg [17:0] R179;
  reg [17:0] R180;
  reg [17:0] R181;
  reg [17:0] R182;
  reg [17:0] R183;
  reg [17:0] R184;
  reg [17:0] R185;
  reg [17:0] R186;
  reg [17:0] R187;
  reg [17:0] R188;
  reg [17:0] R189;
  reg [17:0] R190;
  reg [17:0] R191;
  reg [17:0] R192;
  reg [17:0] R193;
  reg [17:0] R194;
  reg [17:0] R195;
  reg [17:0] R196;
  reg [17:0] R197;
  reg [17:0] R198;
  reg [17:0] R199;
  reg [17:0] R200;
  reg [17:0] R201;
  reg [17:0] R202;
  reg [17:0] R203;
  reg [17:0] R204;
  reg [17:0] R205;
  reg [17:0] R206;
  reg [17:0] R207;
  reg [17:0] R208;
  reg [17:0] R209;
  reg [17:0] R210;
  reg [17:0] R211;
  reg [17:0] R212;
  reg [17:0] R213;
  reg [17:0] R214;
  reg [17:0] R215;
  reg [17:0] R216;
  reg [17:0] R217;
  reg [17:0] R218;
  reg [17:0] R219;
  reg [17:0] R220;
  reg [17:0] R221;
  reg [17:0] R222;
  reg [17:0] R223;
  reg [17:0] R224;
  reg [17:0] R225;
  reg [17:0] R226;
  reg [17:0] R227;
  reg [17:0] R228;
  reg [17:0] R229;
  reg [17:0] R230;
  reg [17:0] R231;
  reg [17:0] R232;
  reg [17:0] R233;
  reg [17:0] R234;
  reg [17:0] R235;
  reg [17:0] R236;
  reg [17:0] R237;
  reg [17:0] R238;
  reg [17:0] R239;
  reg [17:0] R240;
  reg [17:0] R241;
  reg [17:0] R242;
  reg [17:0] R243;
  reg [17:0] R244;
  reg [17:0] R245;
  reg [17:0] R246;
  reg [17:0] R247;
  reg [17:0] R248;
  reg [17:0] R249;
  reg [17:0] R250;
  reg [17:0] R251;
  reg [17:0] R252;
  reg [17:0] R253;
  reg [17:0] R254;
  reg [17:0] R255;
  reg [17:0] R256;
  reg [17:0] R257;
  reg [17:0] R258;
  reg [17:0] R259;
  reg [17:0] R260;
  reg [17:0] R261;
  reg [17:0] R262;
  reg [17:0] R263;
  reg [17:0] R264;
  reg [17:0] R265;
  reg [17:0] R266;
  reg [17:0] R267;
  reg [17:0] R268;
  reg [17:0] R269;
  reg [17:0] R270;
  reg [17:0] R271;
  reg [17:0] R272;
  reg [17:0] R273;
  reg [17:0] R274;
  reg [17:0] R275;
  reg [17:0] R276;
  reg [17:0] R277;
  reg [17:0] R278;
  reg [17:0] R279;
  reg [17:0] R280;
  reg [17:0] R281;
  reg [17:0] R282;
  reg [17:0] R283;
  reg [17:0] R284;
  reg [17:0] R285;
  reg [17:0] R286;
  reg [17:0] R287;
  reg [17:0] R288;
  reg [17:0] R289;
  reg [17:0] R290;
  reg [17:0] R291;
  reg [17:0] R292;
  reg [17:0] R293;
  reg [17:0] R294;
  reg [17:0] R295;
  reg [17:0] R296;
  reg [17:0] R297;
  reg [17:0] R298;
  reg [17:0] R299;
  reg [17:0] R300;
  reg [17:0] R301;
  reg [17:0] R302;
  reg [17:0] R303;
  reg [17:0] R304;
  reg [17:0] R305;
  reg [17:0] R306;
  reg [17:0] R307;
  reg [17:0] R308;
  reg [17:0] R309;
  reg [17:0] R310;
  reg [17:0] R311;
  reg [17:0] R312;
  reg [17:0] R313;
  reg [17:0] R314;
  reg [17:0] R315;
  reg [17:0] R316;
  reg [17:0] R317;
  reg [17:0] R318;
  reg [17:0] R319;
  reg [17:0] R320;
  reg [17:0] R321;
  reg [17:0] R322;
  reg [17:0] R323;
  reg [17:0] R324;
  reg [17:0] R325;
  reg [17:0] R326;
  reg [17:0] R327;
  reg [17:0] R328;
  reg [17:0] R329;
  reg [17:0] R330;
  reg [17:0] R331;
  reg [17:0] R332;
  reg [17:0] R333;
  reg [17:0] R334;
  reg [17:0] R335;
  reg [17:0] R336;
  reg [17:0] R337;
  reg [17:0] R338;
  reg [17:0] R339;
  reg [17:0] R340;
  reg [17:0] R341;
  reg [17:0] R342;
  reg [17:0] R343;
  reg [17:0] R344;
  reg [17:0] R345;
  reg [17:0] R346;
  reg [17:0] R347;
  reg [17:0] R348;
  reg [17:0] R349;
  reg [17:0] R350;
  reg [17:0] R351;
  reg [17:0] R352;
  reg [17:0] R353;
  reg [17:0] R354;
  reg [17:0] R355;
  reg [17:0] R356;
  reg [17:0] R357;
  reg [17:0] R358;
  reg [17:0] R359;
  reg [17:0] R360;
  reg [17:0] R361;
  reg [17:0] R362;
  reg [17:0] R363;
  reg [17:0] R364;
  reg [17:0] R365;
  reg [17:0] R366;
  reg [17:0] R367;
  reg [17:0] R368;
  reg [17:0] R369;
  reg [17:0] R370;
  reg [17:0] R371;
  reg [17:0] R372;
  reg [17:0] R373;
  reg [17:0] R374;
  reg [17:0] R375;
  reg [17:0] R376;
  reg [17:0] R377;
  reg [17:0] R378;
  reg [17:0] R379;
  reg [17:0] R380;
  reg [17:0] R381;
  reg [17:0] R382;
  reg [17:0] R383;
  reg [17:0] R384;
  reg [17:0] R385;
  reg [17:0] R386;
  reg [17:0] R387;
  reg [17:0] R388;
  reg [17:0] R389;
  reg [17:0] R390;
  reg [17:0] R391;
  reg [17:0] R392;
  reg [17:0] R393;
  reg [17:0] R394;
  reg [17:0] R395;
  reg [17:0] R396;
  reg [17:0] R397;
  reg [17:0] R398;
  reg [17:0] R399;
  reg [17:0] R400;
  reg [17:0] R401;
  reg [17:0] R402;
  reg [17:0] R403;
  reg [17:0] R404;
  reg [17:0] R405;
  reg [17:0] R406;
  reg [17:0] R407;
  reg [17:0] R408;
  reg [17:0] R409;
  reg [17:0] R410;
  reg [17:0] R411;
  reg [17:0] R412;
  reg [17:0] R413;
  reg [17:0] R414;
  reg [17:0] R415;
  reg [17:0] R416;
  reg [17:0] R417;
  reg [17:0] R418;
  reg [17:0] R419;
  reg [17:0] R420;
  reg [17:0] R421;
  reg [17:0] R422;
  reg [17:0] R423;
  reg [17:0] R424;
  reg [17:0] R425;
  reg [17:0] R426;
  reg [17:0] R427;
  reg [17:0] R428;
  reg [17:0] R429;
  reg [17:0] R430;
  reg [17:0] R431;
  reg [17:0] R432;
  reg [17:0] R433;
  reg [17:0] R434;
  reg [17:0] R435;
  reg [17:0] R436;
  reg [17:0] R437;
  reg [17:0] R438;
  reg [17:0] R439;
  reg [17:0] R440;
  reg [17:0] R441;
  reg [17:0] R442;
  reg [17:0] R443;
  reg [17:0] R444;
  reg [17:0] R445;
  reg [17:0] R446;
  reg [17:0] R447;
  reg [17:0] R448;
  reg [17:0] R449;
  reg [17:0] R450;
  reg [17:0] R451;
  reg [17:0] R452;
  reg [17:0] R453;
  reg [17:0] R454;
  reg [17:0] R455;
  reg [17:0] R456;
  reg [17:0] R457;
  reg [17:0] R458;
  reg [17:0] R459;
  reg [17:0] R460;
  reg [17:0] R461;
  reg [17:0] R462;
  reg [17:0] R463;
  reg [17:0] R464;
  reg [17:0] R465;
  reg [17:0] R466;
  reg [17:0] R467;
  reg [17:0] R468;
  reg [17:0] R469;
  reg [17:0] R470;
  reg [17:0] zout_0;
  wire[17:0] T471;
  wire[17:0] T472;
  wire[17:0] T473;
  reg [17:0] R474;
  wire[17:0] T475;
  wire[17:0] T1092;
  wire[21:0] T476;
  wire[35:0] T477;
  wire[17:0] T478;
  wire[17:0] T479;
  wire[17:0] T480;
  wire[17:0] T1093;
  wire[21:0] T481;
  wire[35:0] T482;
  wire[17:0] T483;
  wire[17:0] T484;
  wire[17:0] T485;
  wire[17:0] T486;
  wire[17:0] T487;
  reg [17:0] R488;
  wire[17:0] T489;
  wire[17:0] T490;
  reg [17:0] R491;
  reg [17:0] R492;
  reg [17:0] R493;
  reg [17:0] R494;
  reg [17:0] R495;
  reg [17:0] R496;
  reg [17:0] R497;
  reg [17:0] zout_1;
  wire[17:0] T498;
  wire[17:0] T499;
  wire[17:0] T500;
  reg [17:0] R501;
  wire[17:0] T502;
  wire[17:0] T1094;
  wire[21:0] T503;
  wire[35:0] T504;
  wire[17:0] T505;
  wire[17:0] T506;
  wire[17:0] T507;
  wire[17:0] T1095;
  wire[21:0] T508;
  wire[35:0] T509;
  wire[17:0] T510;
  wire[17:0] T511;
  wire[17:0] T512;
  wire[17:0] T513;
  wire[17:0] T514;
  reg [17:0] R515;
  wire[17:0] T516;
  wire[17:0] T517;
  reg [17:0] R518;
  reg [17:0] R519;
  reg [17:0] R520;
  reg [17:0] R521;
  reg [17:0] R522;
  reg [17:0] R523;
  reg [17:0] R524;
  reg [17:0] zout_2;
  wire[17:0] T525;
  wire[17:0] T526;
  wire[17:0] T527;
  reg [17:0] R528;
  wire[17:0] T529;
  wire[17:0] T1096;
  wire[21:0] T530;
  wire[35:0] T531;
  wire[17:0] T532;
  wire[17:0] T533;
  wire[17:0] T534;
  wire[17:0] T1097;
  wire[21:0] T535;
  wire[35:0] T536;
  wire[17:0] T537;
  wire[17:0] T538;
  wire[17:0] T539;
  wire[17:0] T540;
  wire[17:0] T541;
  reg [17:0] R542;
  wire[17:0] T543;
  wire[17:0] T544;
  reg [17:0] R545;
  reg [17:0] R546;
  reg [17:0] R547;
  reg [17:0] R548;
  reg [17:0] R549;
  reg [17:0] R550;
  reg [17:0] R551;
  reg [17:0] yout_0;
  wire[17:0] T552;
  wire[17:0] T553;
  wire[17:0] T554;
  reg [17:0] R555;
  reg [17:0] R556;
  reg [17:0] R557;
  wire[17:0] T558;
  wire[17:0] T1098;
  wire[21:0] T559;
  wire[35:0] T560;
  wire[17:0] T561;
  wire[17:0] T562;
  wire[17:0] T563;
  wire[17:0] T1099;
  wire[21:0] T564;
  wire[35:0] T565;
  wire[17:0] T566;
  wire[17:0] T567;
  wire[17:0] T568;
  wire[17:0] T569;
  wire[17:0] T570;
  reg [17:0] R571;
  reg [17:0] R572;
  reg [17:0] R573;
  reg [17:0] R574;
  reg [17:0] R575;
  reg [17:0] R576;
  reg [17:0] R577;
  reg [17:0] R578;
  wire[17:0] T579;
  reg [17:0] R580;
  reg [17:0] R581;
  reg [17:0] R582;
  reg [17:0] R583;
  reg [17:0] R584;
  wire[17:0] T585;
  reg [17:0] R586;
  reg [17:0] R587;
  reg [17:0] R588;
  reg [17:0] yout_1;
  wire[17:0] T589;
  wire[17:0] T590;
  wire[17:0] T591;
  reg [17:0] R592;
  reg [17:0] R593;
  reg [17:0] R594;
  wire[17:0] T595;
  wire[17:0] T1100;
  wire[21:0] T596;
  wire[35:0] T597;
  wire[17:0] T598;
  wire[17:0] T599;
  wire[17:0] T600;
  wire[17:0] T1101;
  wire[21:0] T601;
  wire[35:0] T602;
  wire[17:0] T603;
  wire[17:0] T604;
  wire[17:0] T605;
  wire[17:0] T606;
  wire[17:0] T607;
  reg [17:0] R608;
  reg [17:0] R609;
  reg [17:0] R610;
  reg [17:0] R611;
  reg [17:0] R612;
  reg [17:0] R613;
  reg [17:0] R614;
  reg [17:0] R615;
  wire[17:0] T616;
  reg [17:0] R617;
  reg [17:0] R618;
  reg [17:0] R619;
  reg [17:0] R620;
  reg [17:0] R621;
  wire[17:0] T622;
  reg [17:0] R623;
  reg [17:0] R624;
  reg [17:0] R625;
  reg [17:0] yout_2;
  wire[17:0] T626;
  wire[17:0] T627;
  wire[17:0] T628;
  reg [17:0] R629;
  reg [17:0] R630;
  reg [17:0] R631;
  wire[17:0] T632;
  wire[17:0] T1102;
  wire[21:0] T633;
  wire[35:0] T634;
  wire[17:0] T635;
  wire[17:0] T636;
  wire[17:0] T637;
  wire[17:0] T1103;
  wire[21:0] T638;
  wire[35:0] T639;
  wire[17:0] T640;
  wire[17:0] T641;
  wire[17:0] T642;
  wire[17:0] T643;
  wire[17:0] T644;
  reg [17:0] R645;
  reg [17:0] R646;
  reg [17:0] R647;
  reg [17:0] R648;
  reg [17:0] R649;
  reg [17:0] R650;
  reg [17:0] R651;
  reg [17:0] R652;
  wire[17:0] T653;
  reg [17:0] R654;
  reg [17:0] R655;
  reg [17:0] R656;
  reg [17:0] R657;
  reg [17:0] R658;
  wire[17:0] T659;
  reg [17:0] R660;
  reg [17:0] R661;
  reg [17:0] R662;
  reg [17:0] yout_3;
  wire[17:0] T663;
  wire[17:0] T664;
  wire[17:0] T665;
  reg [17:0] R666;
  reg [17:0] R667;
  reg [17:0] R668;
  wire[17:0] T669;
  wire[17:0] T1104;
  wire[21:0] T670;
  wire[35:0] T671;
  wire[17:0] T672;
  wire[17:0] T673;
  wire[17:0] T674;
  wire[17:0] T1105;
  wire[21:0] T675;
  wire[35:0] T676;
  wire[17:0] T677;
  wire[17:0] T678;
  wire[17:0] T679;
  wire[17:0] T680;
  wire[17:0] T681;
  reg [17:0] R682;
  reg [17:0] R683;
  reg [17:0] R684;
  reg [17:0] R685;
  reg [17:0] R686;
  reg [17:0] R687;
  reg [17:0] R688;
  reg [17:0] R689;
  wire[17:0] T690;
  reg [17:0] R691;
  reg [17:0] R692;
  reg [17:0] R693;
  reg [17:0] R694;
  reg [17:0] R695;
  wire[17:0] T696;
  reg [17:0] R697;
  reg [17:0] R698;
  reg [17:0] R699;
  reg [17:0] yout_4;
  wire[17:0] T700;
  wire[17:0] T701;
  wire[17:0] T702;
  reg [17:0] R703;
  reg [17:0] R704;
  reg [17:0] R705;
  wire[17:0] T706;
  wire[17:0] T1106;
  wire[21:0] T707;
  wire[35:0] T708;
  wire[17:0] T709;
  wire[17:0] T710;
  wire[17:0] T711;
  wire[17:0] T1107;
  wire[21:0] T712;
  wire[35:0] T713;
  wire[17:0] T714;
  wire[17:0] T715;
  wire[17:0] T716;
  wire[17:0] T717;
  wire[17:0] T718;
  reg [17:0] R719;
  reg [17:0] R720;
  reg [17:0] R721;
  reg [17:0] R722;
  reg [17:0] R723;
  reg [17:0] R724;
  reg [17:0] R725;
  reg [17:0] R726;
  wire[17:0] T727;
  reg [17:0] R728;
  reg [17:0] R729;
  reg [17:0] R730;
  reg [17:0] R731;
  reg [17:0] R732;
  wire[17:0] T733;
  reg [17:0] R734;
  reg [17:0] R735;
  reg [17:0] R736;
  reg [17:0] yout_5;
  wire[17:0] T737;
  wire[17:0] T738;
  wire[17:0] T739;
  reg [17:0] R740;
  reg [17:0] R741;
  reg [17:0] R742;
  wire[17:0] T743;
  wire[17:0] T1108;
  wire[21:0] T744;
  wire[35:0] T745;
  wire[17:0] T746;
  wire[17:0] T747;
  wire[17:0] T748;
  wire[17:0] T1109;
  wire[21:0] T749;
  wire[35:0] T750;
  wire[17:0] T751;
  wire[17:0] T752;
  wire[17:0] T753;
  wire[17:0] T754;
  wire[17:0] T755;
  reg [17:0] R756;
  reg [17:0] R757;
  reg [17:0] R758;
  reg [17:0] R759;
  reg [17:0] R760;
  reg [17:0] R761;
  reg [17:0] R762;
  reg [17:0] R763;
  wire[17:0] T764;
  reg [17:0] R765;
  reg [17:0] R766;
  reg [17:0] R767;
  reg [17:0] R768;
  reg [17:0] R769;
  wire[17:0] T770;
  reg [17:0] R771;
  reg [17:0] R772;
  reg [17:0] R773;
  reg [17:0] yout_6;
  wire[17:0] T774;
  wire[17:0] T775;
  wire[17:0] T776;
  reg [17:0] R777;
  reg [17:0] R778;
  reg [17:0] R779;
  wire[17:0] T780;
  wire[17:0] T1110;
  wire[21:0] T781;
  wire[35:0] T782;
  wire[17:0] T783;
  wire[17:0] T784;
  wire[17:0] T785;
  wire[17:0] T1111;
  wire[21:0] T786;
  wire[35:0] T787;
  wire[17:0] T788;
  wire[17:0] T789;
  wire[17:0] T790;
  wire[17:0] T791;
  wire[17:0] T792;
  reg [17:0] R793;
  reg [17:0] R794;
  reg [17:0] R795;
  reg [17:0] R796;
  reg [17:0] R797;
  reg [17:0] R798;
  reg [17:0] R799;
  reg [17:0] R800;
  wire[17:0] T801;
  reg [17:0] R802;
  reg [17:0] R803;
  reg [17:0] R804;
  reg [17:0] R805;
  reg [17:0] R806;
  wire[17:0] T807;
  reg [17:0] R808;
  reg [17:0] R809;
  reg [17:0] R810;
  reg [17:0] yout_7;
  wire[17:0] T811;
  wire[17:0] T812;
  wire[17:0] T813;
  reg [17:0] R814;
  reg [17:0] R815;
  reg [17:0] R816;
  wire[17:0] T817;
  wire[17:0] T1112;
  wire[21:0] T818;
  wire[35:0] T819;
  wire[17:0] T820;
  wire[17:0] T821;
  wire[17:0] T822;
  wire[17:0] T1113;
  wire[21:0] T823;
  wire[35:0] T824;
  wire[17:0] T825;
  wire[17:0] T826;
  wire[17:0] T827;
  wire[17:0] T828;
  wire[17:0] T829;
  reg [17:0] R830;
  reg [17:0] R831;
  reg [17:0] R832;
  reg [17:0] R833;
  reg [17:0] R834;
  reg [17:0] R835;
  reg [17:0] R836;
  reg [17:0] R837;
  wire[17:0] T838;
  reg [17:0] R839;
  reg [17:0] R840;
  reg [17:0] R841;
  reg [17:0] R842;
  reg [17:0] R843;
  wire[17:0] T844;
  reg [17:0] R845;
  reg [17:0] R846;
  reg [17:0] R847;
  reg [17:0] yout_8;
  wire[17:0] T848;
  wire[17:0] T849;
  wire[17:0] T850;
  reg [17:0] R851;
  reg [17:0] R852;
  reg [17:0] R853;
  wire[17:0] T854;
  wire[17:0] T1114;
  wire[21:0] T855;
  wire[35:0] T856;
  wire[17:0] T857;
  wire[17:0] T858;
  wire[17:0] T859;
  wire[17:0] T1115;
  wire[21:0] T860;
  wire[35:0] T861;
  wire[17:0] T862;
  wire[17:0] T863;
  wire[17:0] T864;
  wire[17:0] T865;
  wire[17:0] T866;
  reg [17:0] R867;
  reg [17:0] R868;
  reg [17:0] R869;
  reg [17:0] R870;
  reg [17:0] R871;
  reg [17:0] R872;
  reg [17:0] R873;
  reg [17:0] R874;
  wire[17:0] T875;
  reg [17:0] R876;
  reg [17:0] R877;
  reg [17:0] R878;
  reg [17:0] R879;
  reg [17:0] R880;
  wire[17:0] T881;
  reg [17:0] R882;
  reg [17:0] R883;
  reg [17:0] R884;
  reg [17:0] yout_9;
  wire[17:0] T885;
  wire[17:0] T886;
  wire[17:0] T887;
  reg [17:0] R888;
  reg [17:0] R889;
  reg [17:0] R890;
  wire[17:0] T891;
  wire[17:0] T1116;
  wire[21:0] T892;
  wire[35:0] T893;
  wire[17:0] T894;
  wire[17:0] T895;
  wire[17:0] T896;
  wire[17:0] T1117;
  wire[21:0] T897;
  wire[35:0] T898;
  wire[17:0] T899;
  wire[17:0] T900;
  wire[17:0] T901;
  wire[17:0] T902;
  wire[17:0] T903;
  reg [17:0] R904;
  reg [17:0] R905;
  reg [17:0] R906;
  reg [17:0] R907;
  reg [17:0] R908;
  reg [17:0] R909;
  reg [17:0] R910;
  reg [17:0] R911;
  wire[17:0] T912;
  reg [17:0] R913;
  reg [17:0] R914;
  reg [17:0] R915;
  reg [17:0] R916;
  reg [17:0] R917;
  wire[17:0] T918;
  reg [17:0] R919;
  reg [17:0] R920;
  reg [17:0] R921;
  reg [17:0] yout_10;
  wire[17:0] T922;
  wire[17:0] T923;
  wire[17:0] T924;
  reg [17:0] R925;
  reg [17:0] R926;
  reg [17:0] R927;
  wire[17:0] T928;
  wire[17:0] T1118;
  wire[21:0] T929;
  wire[35:0] T930;
  wire[17:0] T931;
  wire[17:0] T932;
  wire[17:0] T933;
  wire[17:0] T1119;
  wire[21:0] T934;
  wire[35:0] T935;
  wire[17:0] T936;
  wire[17:0] T937;
  wire[17:0] T938;
  wire[17:0] T939;
  wire[17:0] T940;
  reg [17:0] R941;
  reg [17:0] R942;
  reg [17:0] R943;
  reg [17:0] R944;
  reg [17:0] R945;
  reg [17:0] R946;
  reg [17:0] R947;
  reg [17:0] R948;
  wire[17:0] T949;
  reg [17:0] R950;
  reg [17:0] R951;
  reg [17:0] R952;
  reg [17:0] R953;
  reg [17:0] R954;
  wire[17:0] T955;
  reg [17:0] R956;
  reg [17:0] R957;
  reg [17:0] R958;
  reg [17:0] yout_11;
  wire[17:0] T959;
  wire[17:0] T960;
  wire[17:0] T961;
  reg [17:0] R962;
  reg [17:0] R963;
  reg [17:0] R964;
  wire[17:0] T965;
  wire[17:0] T1120;
  wire[21:0] T966;
  wire[35:0] T967;
  wire[17:0] T968;
  wire[17:0] T969;
  wire[17:0] T970;
  wire[17:0] T1121;
  wire[21:0] T971;
  wire[35:0] T972;
  wire[17:0] T973;
  wire[17:0] T974;
  wire[17:0] T975;
  wire[17:0] T976;
  wire[17:0] T977;
  reg [17:0] R978;
  reg [17:0] R979;
  reg [17:0] R980;
  reg [17:0] R981;
  reg [17:0] R982;
  reg [17:0] R983;
  reg [17:0] R984;
  reg [17:0] R985;
  wire[17:0] T986;
  reg [17:0] R987;
  reg [17:0] R988;
  reg [17:0] R989;
  reg [17:0] R990;
  reg [17:0] R991;
  wire[17:0] T992;
  reg [17:0] R993;
  reg [17:0] R994;
  reg [17:0] R995;
  reg [17:0] xout_0;
  wire[17:0] T996;
  wire[17:0] T997;
  wire[17:0] T998;
  reg [17:0] R999;
  reg [17:0] R1000;
  reg [17:0] R1001;
  wire[17:0] T1002;
  wire[17:0] T1122;
  wire[21:0] T1003;
  wire[35:0] T1004;
  wire[17:0] T1005;
  wire[17:0] T1006;
  wire[17:0] T1007;
  wire[17:0] T1008;
  wire[17:0] T1009;
  reg [17:0] R1010;
  reg [17:0] R1011;
  reg [17:0] R1012;
  reg [17:0] R1013;
  reg [17:0] R1014;
  reg [17:0] R1015;
  reg [17:0] R1016;
  reg [17:0] R1017;
  reg [17:0] R1018;
  reg [17:0] R1019;
  reg [17:0] R1020;
  reg [17:0] R1021;
  reg [17:0] R1022;
  wire[17:0] T1023;
  wire[17:0] T1024;
  reg [17:0] R1025;
  reg [17:0] R1026;
  reg [17:0] R1027;
  reg [17:0] xout_1;
  wire[17:0] T1028;
  wire[17:0] T1029;
  wire[17:0] T1030;
  reg [17:0] R1031;
  reg [17:0] R1032;
  reg [17:0] R1033;
  wire[17:0] T1034;
  wire[17:0] T1123;
  wire[21:0] T1035;
  wire[35:0] T1036;
  wire[17:0] T1037;
  wire[17:0] T1038;
  wire[17:0] T1039;
  wire[17:0] T1040;
  wire[17:0] T1041;
  reg [17:0] R1042;
  reg [17:0] R1043;
  reg [17:0] R1044;
  reg [17:0] R1045;
  reg [17:0] R1046;
  reg [17:0] R1047;
  reg [17:0] R1048;
  reg [17:0] R1049;
  reg [17:0] R1050;
  reg [17:0] R1051;
  reg [17:0] R1052;
  reg [17:0] R1053;
  reg [17:0] R1054;
  wire[17:0] T1055;
  wire[17:0] T1056;
  reg [17:0] R1057;
  reg [17:0] R1058;
  reg [17:0] R1059;
  reg [17:0] xout_2;
  wire[17:0] T1060;
  wire[17:0] T1061;
  wire[17:0] T1062;
  reg [17:0] R1063;
  reg [17:0] R1064;
  reg [17:0] R1065;
  wire[17:0] T1066;
  wire[17:0] T1124;
  wire[21:0] T1067;
  wire[35:0] T1068;
  wire[17:0] T1069;
  wire[17:0] T1070;
  wire[17:0] T1071;
  wire[17:0] T1072;
  wire[17:0] T1073;
  reg [17:0] R1074;
  reg [17:0] R1075;
  reg [17:0] R1076;
  reg [17:0] R1077;
  reg [17:0] R1078;
  reg [17:0] R1079;
  reg [17:0] R1080;
  reg [17:0] R1081;
  reg [17:0] R1082;
  reg [17:0] R1083;
  reg [17:0] R1084;
  reg [17:0] R1085;
  reg [17:0] R1086;
  wire[17:0] T1087;
  wire[17:0] T1088;
  reg [17:0] R1089;
  reg [17:0] R1090;
  reg [17:0] R1091;
  wire[17:0] MatrixVectorMultModule_io_o_2;
  wire[17:0] MatrixVectorMultModule_io_o_1;
  wire[17:0] MatrixVectorMultModule_io_o_0;
  wire[17:0] XNetModule_io_o_2;
  wire[17:0] XNetModule_io_o_1;
  wire[17:0] XNetModule_io_o_0;
  wire[17:0] YNetModule_io_o_11;
  wire[17:0] YNetModule_io_o_10;
  wire[17:0] YNetModule_io_o_9;
  wire[17:0] YNetModule_io_o_8;
  wire[17:0] YNetModule_io_o_7;
  wire[17:0] YNetModule_io_o_6;
  wire[17:0] YNetModule_io_o_5;
  wire[17:0] YNetModule_io_o_4;
  wire[17:0] YNetModule_io_o_3;
  wire[17:0] YNetModule_io_o_2;
  wire[17:0] YNetModule_io_o_1;
  wire[17:0] YNetModule_io_o_0;
  wire[17:0] ZNetModule_io_o_2;
  wire[17:0] ZNetModule_io_o_1;
  wire[17:0] ZNetModule_io_o_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
    R2 = {1{$random}};
    R3 = {1{$random}};
    R4 = {1{$random}};
    R5 = {1{$random}};
    R6 = {1{$random}};
    R7 = {1{$random}};
    R8 = {1{$random}};
    R9 = {1{$random}};
    R10 = {1{$random}};
    R11 = {1{$random}};
    R12 = {1{$random}};
    R13 = {1{$random}};
    R14 = {1{$random}};
    R15 = {1{$random}};
    R16 = {1{$random}};
    R17 = {1{$random}};
    R18 = {1{$random}};
    R19 = {1{$random}};
    R20 = {1{$random}};
    R21 = {1{$random}};
    R22 = {1{$random}};
    R23 = {1{$random}};
    R24 = {1{$random}};
    R25 = {1{$random}};
    R26 = {1{$random}};
    R27 = {1{$random}};
    R28 = {1{$random}};
    R29 = {1{$random}};
    R30 = {1{$random}};
    R31 = {1{$random}};
    R32 = {1{$random}};
    R33 = {1{$random}};
    R34 = {1{$random}};
    R35 = {1{$random}};
    R36 = {1{$random}};
    R37 = {1{$random}};
    R38 = {1{$random}};
    R39 = {1{$random}};
    R40 = {1{$random}};
    R41 = {1{$random}};
    R42 = {1{$random}};
    R43 = {1{$random}};
    R44 = {1{$random}};
    R45 = {1{$random}};
    R46 = {1{$random}};
    R47 = {1{$random}};
    R48 = {1{$random}};
    R49 = {1{$random}};
    R50 = {1{$random}};
    R51 = {1{$random}};
    R52 = {1{$random}};
    R53 = {1{$random}};
    R54 = {1{$random}};
    R55 = {1{$random}};
    R56 = {1{$random}};
    R57 = {1{$random}};
    R58 = {1{$random}};
    R59 = {1{$random}};
    R60 = {1{$random}};
    R61 = {1{$random}};
    R62 = {1{$random}};
    R63 = {1{$random}};
    R64 = {1{$random}};
    R65 = {1{$random}};
    R66 = {1{$random}};
    R67 = {1{$random}};
    R68 = {1{$random}};
    R69 = {1{$random}};
    R70 = {1{$random}};
    R71 = {1{$random}};
    R72 = {1{$random}};
    R73 = {1{$random}};
    R74 = {1{$random}};
    R75 = {1{$random}};
    R76 = {1{$random}};
    R77 = {1{$random}};
    R78 = {1{$random}};
    R79 = {1{$random}};
    R80 = {1{$random}};
    R81 = {1{$random}};
    R82 = {1{$random}};
    R83 = {1{$random}};
    R84 = {1{$random}};
    R85 = {1{$random}};
    R86 = {1{$random}};
    R87 = {1{$random}};
    R88 = {1{$random}};
    R89 = {1{$random}};
    R90 = {1{$random}};
    R91 = {1{$random}};
    R92 = {1{$random}};
    R93 = {1{$random}};
    R94 = {1{$random}};
    R95 = {1{$random}};
    R96 = {1{$random}};
    R97 = {1{$random}};
    R98 = {1{$random}};
    R99 = {1{$random}};
    R100 = {1{$random}};
    R101 = {1{$random}};
    R102 = {1{$random}};
    R103 = {1{$random}};
    R104 = {1{$random}};
    R105 = {1{$random}};
    R106 = {1{$random}};
    R107 = {1{$random}};
    R108 = {1{$random}};
    R109 = {1{$random}};
    R110 = {1{$random}};
    R111 = {1{$random}};
    R112 = {1{$random}};
    R113 = {1{$random}};
    R114 = {1{$random}};
    R115 = {1{$random}};
    R116 = {1{$random}};
    R117 = {1{$random}};
    R118 = {1{$random}};
    R119 = {1{$random}};
    R120 = {1{$random}};
    R121 = {1{$random}};
    R122 = {1{$random}};
    R123 = {1{$random}};
    R124 = {1{$random}};
    R125 = {1{$random}};
    R126 = {1{$random}};
    R127 = {1{$random}};
    R128 = {1{$random}};
    R129 = {1{$random}};
    R130 = {1{$random}};
    R131 = {1{$random}};
    R132 = {1{$random}};
    R133 = {1{$random}};
    R134 = {1{$random}};
    R135 = {1{$random}};
    R136 = {1{$random}};
    R137 = {1{$random}};
    R138 = {1{$random}};
    R139 = {1{$random}};
    R140 = {1{$random}};
    R141 = {1{$random}};
    R142 = {1{$random}};
    R143 = {1{$random}};
    R144 = {1{$random}};
    R145 = {1{$random}};
    R146 = {1{$random}};
    R147 = {1{$random}};
    R148 = {1{$random}};
    R149 = {1{$random}};
    R150 = {1{$random}};
    R151 = {1{$random}};
    R152 = {1{$random}};
    R153 = {1{$random}};
    R154 = {1{$random}};
    R155 = {1{$random}};
    R156 = {1{$random}};
    R157 = {1{$random}};
    R158 = {1{$random}};
    R159 = {1{$random}};
    R160 = {1{$random}};
    R161 = {1{$random}};
    R162 = {1{$random}};
    R163 = {1{$random}};
    R164 = {1{$random}};
    R165 = {1{$random}};
    R166 = {1{$random}};
    R167 = {1{$random}};
    R168 = {1{$random}};
    R169 = {1{$random}};
    R170 = {1{$random}};
    R171 = {1{$random}};
    R172 = {1{$random}};
    R173 = {1{$random}};
    R174 = {1{$random}};
    R175 = {1{$random}};
    R176 = {1{$random}};
    R177 = {1{$random}};
    R178 = {1{$random}};
    R179 = {1{$random}};
    R180 = {1{$random}};
    R181 = {1{$random}};
    R182 = {1{$random}};
    R183 = {1{$random}};
    R184 = {1{$random}};
    R185 = {1{$random}};
    R186 = {1{$random}};
    R187 = {1{$random}};
    R188 = {1{$random}};
    R189 = {1{$random}};
    R190 = {1{$random}};
    R191 = {1{$random}};
    R192 = {1{$random}};
    R193 = {1{$random}};
    R194 = {1{$random}};
    R195 = {1{$random}};
    R196 = {1{$random}};
    R197 = {1{$random}};
    R198 = {1{$random}};
    R199 = {1{$random}};
    R200 = {1{$random}};
    R201 = {1{$random}};
    R202 = {1{$random}};
    R203 = {1{$random}};
    R204 = {1{$random}};
    R205 = {1{$random}};
    R206 = {1{$random}};
    R207 = {1{$random}};
    R208 = {1{$random}};
    R209 = {1{$random}};
    R210 = {1{$random}};
    R211 = {1{$random}};
    R212 = {1{$random}};
    R213 = {1{$random}};
    R214 = {1{$random}};
    R215 = {1{$random}};
    R216 = {1{$random}};
    R217 = {1{$random}};
    R218 = {1{$random}};
    R219 = {1{$random}};
    R220 = {1{$random}};
    R221 = {1{$random}};
    R222 = {1{$random}};
    R223 = {1{$random}};
    R224 = {1{$random}};
    R225 = {1{$random}};
    R226 = {1{$random}};
    R227 = {1{$random}};
    R228 = {1{$random}};
    R229 = {1{$random}};
    R230 = {1{$random}};
    R231 = {1{$random}};
    R232 = {1{$random}};
    R233 = {1{$random}};
    R234 = {1{$random}};
    R235 = {1{$random}};
    R236 = {1{$random}};
    R237 = {1{$random}};
    R238 = {1{$random}};
    R239 = {1{$random}};
    R240 = {1{$random}};
    R241 = {1{$random}};
    R242 = {1{$random}};
    R243 = {1{$random}};
    R244 = {1{$random}};
    R245 = {1{$random}};
    R246 = {1{$random}};
    R247 = {1{$random}};
    R248 = {1{$random}};
    R249 = {1{$random}};
    R250 = {1{$random}};
    R251 = {1{$random}};
    R252 = {1{$random}};
    R253 = {1{$random}};
    R254 = {1{$random}};
    R255 = {1{$random}};
    R256 = {1{$random}};
    R257 = {1{$random}};
    R258 = {1{$random}};
    R259 = {1{$random}};
    R260 = {1{$random}};
    R261 = {1{$random}};
    R262 = {1{$random}};
    R263 = {1{$random}};
    R264 = {1{$random}};
    R265 = {1{$random}};
    R266 = {1{$random}};
    R267 = {1{$random}};
    R268 = {1{$random}};
    R269 = {1{$random}};
    R270 = {1{$random}};
    R271 = {1{$random}};
    R272 = {1{$random}};
    R273 = {1{$random}};
    R274 = {1{$random}};
    R275 = {1{$random}};
    R276 = {1{$random}};
    R277 = {1{$random}};
    R278 = {1{$random}};
    R279 = {1{$random}};
    R280 = {1{$random}};
    R281 = {1{$random}};
    R282 = {1{$random}};
    R283 = {1{$random}};
    R284 = {1{$random}};
    R285 = {1{$random}};
    R286 = {1{$random}};
    R287 = {1{$random}};
    R288 = {1{$random}};
    R289 = {1{$random}};
    R290 = {1{$random}};
    R291 = {1{$random}};
    R292 = {1{$random}};
    R293 = {1{$random}};
    R294 = {1{$random}};
    R295 = {1{$random}};
    R296 = {1{$random}};
    R297 = {1{$random}};
    R298 = {1{$random}};
    R299 = {1{$random}};
    R300 = {1{$random}};
    R301 = {1{$random}};
    R302 = {1{$random}};
    R303 = {1{$random}};
    R304 = {1{$random}};
    R305 = {1{$random}};
    R306 = {1{$random}};
    R307 = {1{$random}};
    R308 = {1{$random}};
    R309 = {1{$random}};
    R310 = {1{$random}};
    R311 = {1{$random}};
    R312 = {1{$random}};
    R313 = {1{$random}};
    R314 = {1{$random}};
    R315 = {1{$random}};
    R316 = {1{$random}};
    R317 = {1{$random}};
    R318 = {1{$random}};
    R319 = {1{$random}};
    R320 = {1{$random}};
    R321 = {1{$random}};
    R322 = {1{$random}};
    R323 = {1{$random}};
    R324 = {1{$random}};
    R325 = {1{$random}};
    R326 = {1{$random}};
    R327 = {1{$random}};
    R328 = {1{$random}};
    R329 = {1{$random}};
    R330 = {1{$random}};
    R331 = {1{$random}};
    R332 = {1{$random}};
    R333 = {1{$random}};
    R334 = {1{$random}};
    R335 = {1{$random}};
    R336 = {1{$random}};
    R337 = {1{$random}};
    R338 = {1{$random}};
    R339 = {1{$random}};
    R340 = {1{$random}};
    R341 = {1{$random}};
    R342 = {1{$random}};
    R343 = {1{$random}};
    R344 = {1{$random}};
    R345 = {1{$random}};
    R346 = {1{$random}};
    R347 = {1{$random}};
    R348 = {1{$random}};
    R349 = {1{$random}};
    R350 = {1{$random}};
    R351 = {1{$random}};
    R352 = {1{$random}};
    R353 = {1{$random}};
    R354 = {1{$random}};
    R355 = {1{$random}};
    R356 = {1{$random}};
    R357 = {1{$random}};
    R358 = {1{$random}};
    R359 = {1{$random}};
    R360 = {1{$random}};
    R361 = {1{$random}};
    R362 = {1{$random}};
    R363 = {1{$random}};
    R364 = {1{$random}};
    R365 = {1{$random}};
    R366 = {1{$random}};
    R367 = {1{$random}};
    R368 = {1{$random}};
    R369 = {1{$random}};
    R370 = {1{$random}};
    R371 = {1{$random}};
    R372 = {1{$random}};
    R373 = {1{$random}};
    R374 = {1{$random}};
    R375 = {1{$random}};
    R376 = {1{$random}};
    R377 = {1{$random}};
    R378 = {1{$random}};
    R379 = {1{$random}};
    R380 = {1{$random}};
    R381 = {1{$random}};
    R382 = {1{$random}};
    R383 = {1{$random}};
    R384 = {1{$random}};
    R385 = {1{$random}};
    R386 = {1{$random}};
    R387 = {1{$random}};
    R388 = {1{$random}};
    R389 = {1{$random}};
    R390 = {1{$random}};
    R391 = {1{$random}};
    R392 = {1{$random}};
    R393 = {1{$random}};
    R394 = {1{$random}};
    R395 = {1{$random}};
    R396 = {1{$random}};
    R397 = {1{$random}};
    R398 = {1{$random}};
    R399 = {1{$random}};
    R400 = {1{$random}};
    R401 = {1{$random}};
    R402 = {1{$random}};
    R403 = {1{$random}};
    R404 = {1{$random}};
    R405 = {1{$random}};
    R406 = {1{$random}};
    R407 = {1{$random}};
    R408 = {1{$random}};
    R409 = {1{$random}};
    R410 = {1{$random}};
    R411 = {1{$random}};
    R412 = {1{$random}};
    R413 = {1{$random}};
    R414 = {1{$random}};
    R415 = {1{$random}};
    R416 = {1{$random}};
    R417 = {1{$random}};
    R418 = {1{$random}};
    R419 = {1{$random}};
    R420 = {1{$random}};
    R421 = {1{$random}};
    R422 = {1{$random}};
    R423 = {1{$random}};
    R424 = {1{$random}};
    R425 = {1{$random}};
    R426 = {1{$random}};
    R427 = {1{$random}};
    R428 = {1{$random}};
    R429 = {1{$random}};
    R430 = {1{$random}};
    R431 = {1{$random}};
    R432 = {1{$random}};
    R433 = {1{$random}};
    R434 = {1{$random}};
    R435 = {1{$random}};
    R436 = {1{$random}};
    R437 = {1{$random}};
    R438 = {1{$random}};
    R439 = {1{$random}};
    R440 = {1{$random}};
    R441 = {1{$random}};
    R442 = {1{$random}};
    R443 = {1{$random}};
    R444 = {1{$random}};
    R445 = {1{$random}};
    R446 = {1{$random}};
    R447 = {1{$random}};
    R448 = {1{$random}};
    R449 = {1{$random}};
    R450 = {1{$random}};
    R451 = {1{$random}};
    R452 = {1{$random}};
    R453 = {1{$random}};
    R454 = {1{$random}};
    R455 = {1{$random}};
    R456 = {1{$random}};
    R457 = {1{$random}};
    R458 = {1{$random}};
    R459 = {1{$random}};
    R460 = {1{$random}};
    R461 = {1{$random}};
    R462 = {1{$random}};
    R463 = {1{$random}};
    R464 = {1{$random}};
    R465 = {1{$random}};
    R466 = {1{$random}};
    R467 = {1{$random}};
    R468 = {1{$random}};
    R469 = {1{$random}};
    R470 = {1{$random}};
    zout_0 = {1{$random}};
    R474 = {1{$random}};
    R488 = {1{$random}};
    R491 = {1{$random}};
    R492 = {1{$random}};
    R493 = {1{$random}};
    R494 = {1{$random}};
    R495 = {1{$random}};
    R496 = {1{$random}};
    R497 = {1{$random}};
    zout_1 = {1{$random}};
    R501 = {1{$random}};
    R515 = {1{$random}};
    R518 = {1{$random}};
    R519 = {1{$random}};
    R520 = {1{$random}};
    R521 = {1{$random}};
    R522 = {1{$random}};
    R523 = {1{$random}};
    R524 = {1{$random}};
    zout_2 = {1{$random}};
    R528 = {1{$random}};
    R542 = {1{$random}};
    R545 = {1{$random}};
    R546 = {1{$random}};
    R547 = {1{$random}};
    R548 = {1{$random}};
    R549 = {1{$random}};
    R550 = {1{$random}};
    R551 = {1{$random}};
    yout_0 = {1{$random}};
    R555 = {1{$random}};
    R556 = {1{$random}};
    R557 = {1{$random}};
    R571 = {1{$random}};
    R572 = {1{$random}};
    R573 = {1{$random}};
    R574 = {1{$random}};
    R575 = {1{$random}};
    R576 = {1{$random}};
    R577 = {1{$random}};
    R578 = {1{$random}};
    R580 = {1{$random}};
    R581 = {1{$random}};
    R582 = {1{$random}};
    R583 = {1{$random}};
    R584 = {1{$random}};
    R586 = {1{$random}};
    R587 = {1{$random}};
    R588 = {1{$random}};
    yout_1 = {1{$random}};
    R592 = {1{$random}};
    R593 = {1{$random}};
    R594 = {1{$random}};
    R608 = {1{$random}};
    R609 = {1{$random}};
    R610 = {1{$random}};
    R611 = {1{$random}};
    R612 = {1{$random}};
    R613 = {1{$random}};
    R614 = {1{$random}};
    R615 = {1{$random}};
    R617 = {1{$random}};
    R618 = {1{$random}};
    R619 = {1{$random}};
    R620 = {1{$random}};
    R621 = {1{$random}};
    R623 = {1{$random}};
    R624 = {1{$random}};
    R625 = {1{$random}};
    yout_2 = {1{$random}};
    R629 = {1{$random}};
    R630 = {1{$random}};
    R631 = {1{$random}};
    R645 = {1{$random}};
    R646 = {1{$random}};
    R647 = {1{$random}};
    R648 = {1{$random}};
    R649 = {1{$random}};
    R650 = {1{$random}};
    R651 = {1{$random}};
    R652 = {1{$random}};
    R654 = {1{$random}};
    R655 = {1{$random}};
    R656 = {1{$random}};
    R657 = {1{$random}};
    R658 = {1{$random}};
    R660 = {1{$random}};
    R661 = {1{$random}};
    R662 = {1{$random}};
    yout_3 = {1{$random}};
    R666 = {1{$random}};
    R667 = {1{$random}};
    R668 = {1{$random}};
    R682 = {1{$random}};
    R683 = {1{$random}};
    R684 = {1{$random}};
    R685 = {1{$random}};
    R686 = {1{$random}};
    R687 = {1{$random}};
    R688 = {1{$random}};
    R689 = {1{$random}};
    R691 = {1{$random}};
    R692 = {1{$random}};
    R693 = {1{$random}};
    R694 = {1{$random}};
    R695 = {1{$random}};
    R697 = {1{$random}};
    R698 = {1{$random}};
    R699 = {1{$random}};
    yout_4 = {1{$random}};
    R703 = {1{$random}};
    R704 = {1{$random}};
    R705 = {1{$random}};
    R719 = {1{$random}};
    R720 = {1{$random}};
    R721 = {1{$random}};
    R722 = {1{$random}};
    R723 = {1{$random}};
    R724 = {1{$random}};
    R725 = {1{$random}};
    R726 = {1{$random}};
    R728 = {1{$random}};
    R729 = {1{$random}};
    R730 = {1{$random}};
    R731 = {1{$random}};
    R732 = {1{$random}};
    R734 = {1{$random}};
    R735 = {1{$random}};
    R736 = {1{$random}};
    yout_5 = {1{$random}};
    R740 = {1{$random}};
    R741 = {1{$random}};
    R742 = {1{$random}};
    R756 = {1{$random}};
    R757 = {1{$random}};
    R758 = {1{$random}};
    R759 = {1{$random}};
    R760 = {1{$random}};
    R761 = {1{$random}};
    R762 = {1{$random}};
    R763 = {1{$random}};
    R765 = {1{$random}};
    R766 = {1{$random}};
    R767 = {1{$random}};
    R768 = {1{$random}};
    R769 = {1{$random}};
    R771 = {1{$random}};
    R772 = {1{$random}};
    R773 = {1{$random}};
    yout_6 = {1{$random}};
    R777 = {1{$random}};
    R778 = {1{$random}};
    R779 = {1{$random}};
    R793 = {1{$random}};
    R794 = {1{$random}};
    R795 = {1{$random}};
    R796 = {1{$random}};
    R797 = {1{$random}};
    R798 = {1{$random}};
    R799 = {1{$random}};
    R800 = {1{$random}};
    R802 = {1{$random}};
    R803 = {1{$random}};
    R804 = {1{$random}};
    R805 = {1{$random}};
    R806 = {1{$random}};
    R808 = {1{$random}};
    R809 = {1{$random}};
    R810 = {1{$random}};
    yout_7 = {1{$random}};
    R814 = {1{$random}};
    R815 = {1{$random}};
    R816 = {1{$random}};
    R830 = {1{$random}};
    R831 = {1{$random}};
    R832 = {1{$random}};
    R833 = {1{$random}};
    R834 = {1{$random}};
    R835 = {1{$random}};
    R836 = {1{$random}};
    R837 = {1{$random}};
    R839 = {1{$random}};
    R840 = {1{$random}};
    R841 = {1{$random}};
    R842 = {1{$random}};
    R843 = {1{$random}};
    R845 = {1{$random}};
    R846 = {1{$random}};
    R847 = {1{$random}};
    yout_8 = {1{$random}};
    R851 = {1{$random}};
    R852 = {1{$random}};
    R853 = {1{$random}};
    R867 = {1{$random}};
    R868 = {1{$random}};
    R869 = {1{$random}};
    R870 = {1{$random}};
    R871 = {1{$random}};
    R872 = {1{$random}};
    R873 = {1{$random}};
    R874 = {1{$random}};
    R876 = {1{$random}};
    R877 = {1{$random}};
    R878 = {1{$random}};
    R879 = {1{$random}};
    R880 = {1{$random}};
    R882 = {1{$random}};
    R883 = {1{$random}};
    R884 = {1{$random}};
    yout_9 = {1{$random}};
    R888 = {1{$random}};
    R889 = {1{$random}};
    R890 = {1{$random}};
    R904 = {1{$random}};
    R905 = {1{$random}};
    R906 = {1{$random}};
    R907 = {1{$random}};
    R908 = {1{$random}};
    R909 = {1{$random}};
    R910 = {1{$random}};
    R911 = {1{$random}};
    R913 = {1{$random}};
    R914 = {1{$random}};
    R915 = {1{$random}};
    R916 = {1{$random}};
    R917 = {1{$random}};
    R919 = {1{$random}};
    R920 = {1{$random}};
    R921 = {1{$random}};
    yout_10 = {1{$random}};
    R925 = {1{$random}};
    R926 = {1{$random}};
    R927 = {1{$random}};
    R941 = {1{$random}};
    R942 = {1{$random}};
    R943 = {1{$random}};
    R944 = {1{$random}};
    R945 = {1{$random}};
    R946 = {1{$random}};
    R947 = {1{$random}};
    R948 = {1{$random}};
    R950 = {1{$random}};
    R951 = {1{$random}};
    R952 = {1{$random}};
    R953 = {1{$random}};
    R954 = {1{$random}};
    R956 = {1{$random}};
    R957 = {1{$random}};
    R958 = {1{$random}};
    yout_11 = {1{$random}};
    R962 = {1{$random}};
    R963 = {1{$random}};
    R964 = {1{$random}};
    R978 = {1{$random}};
    R979 = {1{$random}};
    R980 = {1{$random}};
    R981 = {1{$random}};
    R982 = {1{$random}};
    R983 = {1{$random}};
    R984 = {1{$random}};
    R985 = {1{$random}};
    R987 = {1{$random}};
    R988 = {1{$random}};
    R989 = {1{$random}};
    R990 = {1{$random}};
    R991 = {1{$random}};
    R993 = {1{$random}};
    R994 = {1{$random}};
    R995 = {1{$random}};
    xout_0 = {1{$random}};
    R999 = {1{$random}};
    R1000 = {1{$random}};
    R1001 = {1{$random}};
    R1010 = {1{$random}};
    R1011 = {1{$random}};
    R1012 = {1{$random}};
    R1013 = {1{$random}};
    R1014 = {1{$random}};
    R1015 = {1{$random}};
    R1016 = {1{$random}};
    R1017 = {1{$random}};
    R1018 = {1{$random}};
    R1019 = {1{$random}};
    R1020 = {1{$random}};
    R1021 = {1{$random}};
    R1022 = {1{$random}};
    R1025 = {1{$random}};
    R1026 = {1{$random}};
    R1027 = {1{$random}};
    xout_1 = {1{$random}};
    R1031 = {1{$random}};
    R1032 = {1{$random}};
    R1033 = {1{$random}};
    R1042 = {1{$random}};
    R1043 = {1{$random}};
    R1044 = {1{$random}};
    R1045 = {1{$random}};
    R1046 = {1{$random}};
    R1047 = {1{$random}};
    R1048 = {1{$random}};
    R1049 = {1{$random}};
    R1050 = {1{$random}};
    R1051 = {1{$random}};
    R1052 = {1{$random}};
    R1053 = {1{$random}};
    R1054 = {1{$random}};
    R1057 = {1{$random}};
    R1058 = {1{$random}};
    R1059 = {1{$random}};
    xout_2 = {1{$random}};
    R1063 = {1{$random}};
    R1064 = {1{$random}};
    R1065 = {1{$random}};
    R1074 = {1{$random}};
    R1075 = {1{$random}};
    R1076 = {1{$random}};
    R1077 = {1{$random}};
    R1078 = {1{$random}};
    R1079 = {1{$random}};
    R1080 = {1{$random}};
    R1081 = {1{$random}};
    R1082 = {1{$random}};
    R1083 = {1{$random}};
    R1084 = {1{$random}};
    R1085 = {1{$random}};
    R1086 = {1{$random}};
    R1089 = {1{$random}};
    R1090 = {1{$random}};
    R1091 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_zout_0 = zout_0;
  assign T471 = T472;
  assign T472 = T490 + T473;
  assign T473 = R474;
  assign T475 = T1092;
  assign T1092 = T476[5'h11:1'h0];
  assign T476 = $signed(T477) >>> 4'he;
  assign T477 = $signed(T479) * $signed(T478);
  assign T478 = 18'h8000;
  assign T479 = T480;
  assign T480 = T1093;
  assign T1093 = T481[5'h11:1'h0];
  assign T481 = $signed(T482) >>> 4'he;
  assign T482 = $signed(T484) * $signed(T483);
  assign T483 = io_lbda;
  assign T484 = T485;
  assign T485 = T486;
  assign T486 = T489 - T487;
  assign T487 = R488;
  assign T489 = MatrixVectorMultModule_io_o_0;
  assign T490 = R491;
  assign io_zout_1 = zout_1;
  assign T498 = T499;
  assign T499 = T517 + T500;
  assign T500 = R501;
  assign T502 = T1094;
  assign T1094 = T503[5'h11:1'h0];
  assign T503 = $signed(T504) >>> 4'he;
  assign T504 = $signed(T506) * $signed(T505);
  assign T505 = 18'h8000;
  assign T506 = T507;
  assign T507 = T1095;
  assign T1095 = T508[5'h11:1'h0];
  assign T508 = $signed(T509) >>> 4'he;
  assign T509 = $signed(T511) * $signed(T510);
  assign T510 = io_lbda;
  assign T511 = T512;
  assign T512 = T513;
  assign T513 = T516 - T514;
  assign T514 = R515;
  assign T516 = MatrixVectorMultModule_io_o_1;
  assign T517 = R518;
  assign io_zout_2 = zout_2;
  assign T525 = T526;
  assign T526 = T544 + T527;
  assign T527 = R528;
  assign T529 = T1096;
  assign T1096 = T530[5'h11:1'h0];
  assign T530 = $signed(T531) >>> 4'he;
  assign T531 = $signed(T533) * $signed(T532);
  assign T532 = 18'h8000;
  assign T533 = T534;
  assign T534 = T1097;
  assign T1097 = T535[5'h11:1'h0];
  assign T535 = $signed(T536) >>> 4'he;
  assign T536 = $signed(T538) * $signed(T537);
  assign T537 = io_lbda;
  assign T538 = T539;
  assign T539 = T540;
  assign T540 = T543 - T541;
  assign T541 = R542;
  assign T543 = MatrixVectorMultModule_io_o_2;
  assign T544 = R545;
  assign io_yout_0 = yout_0;
  assign T552 = T553;
  assign T553 = T585 + T554;
  assign T554 = R555;
  assign T558 = T1098;
  assign T1098 = T559[5'h11:1'h0];
  assign T559 = $signed(T560) >>> 4'he;
  assign T560 = $signed(T562) * $signed(T561);
  assign T561 = 18'h8000;
  assign T562 = T563;
  assign T563 = T1099;
  assign T1099 = T564[5'h11:1'h0];
  assign T564 = $signed(T565) >>> 4'he;
  assign T565 = $signed(T567) * $signed(T566);
  assign T566 = io_lbda;
  assign T567 = T568;
  assign T568 = T569;
  assign T569 = T579 - T570;
  assign T570 = R571;
  assign T579 = R580;
  assign T585 = R586;
  assign io_yout_1 = yout_1;
  assign T589 = T590;
  assign T590 = T622 + T591;
  assign T591 = R592;
  assign T595 = T1100;
  assign T1100 = T596[5'h11:1'h0];
  assign T596 = $signed(T597) >>> 4'he;
  assign T597 = $signed(T599) * $signed(T598);
  assign T598 = 18'h8000;
  assign T599 = T600;
  assign T600 = T1101;
  assign T1101 = T601[5'h11:1'h0];
  assign T601 = $signed(T602) >>> 4'he;
  assign T602 = $signed(T604) * $signed(T603);
  assign T603 = io_lbda;
  assign T604 = T605;
  assign T605 = T606;
  assign T606 = T616 - T607;
  assign T607 = R608;
  assign T616 = R617;
  assign T622 = R623;
  assign io_yout_2 = yout_2;
  assign T626 = T627;
  assign T627 = T659 + T628;
  assign T628 = R629;
  assign T632 = T1102;
  assign T1102 = T633[5'h11:1'h0];
  assign T633 = $signed(T634) >>> 4'he;
  assign T634 = $signed(T636) * $signed(T635);
  assign T635 = 18'h8000;
  assign T636 = T637;
  assign T637 = T1103;
  assign T1103 = T638[5'h11:1'h0];
  assign T638 = $signed(T639) >>> 4'he;
  assign T639 = $signed(T641) * $signed(T640);
  assign T640 = io_lbda;
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = T653 - T644;
  assign T644 = R645;
  assign T653 = R654;
  assign T659 = R660;
  assign io_yout_3 = yout_3;
  assign T663 = T664;
  assign T664 = T696 + T665;
  assign T665 = R666;
  assign T669 = T1104;
  assign T1104 = T670[5'h11:1'h0];
  assign T670 = $signed(T671) >>> 4'he;
  assign T671 = $signed(T673) * $signed(T672);
  assign T672 = 18'h8000;
  assign T673 = T674;
  assign T674 = T1105;
  assign T1105 = T675[5'h11:1'h0];
  assign T675 = $signed(T676) >>> 4'he;
  assign T676 = $signed(T678) * $signed(T677);
  assign T677 = io_lbda;
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T690 - T681;
  assign T681 = R682;
  assign T690 = R691;
  assign T696 = R697;
  assign io_yout_4 = yout_4;
  assign T700 = T701;
  assign T701 = T733 + T702;
  assign T702 = R703;
  assign T706 = T1106;
  assign T1106 = T707[5'h11:1'h0];
  assign T707 = $signed(T708) >>> 4'he;
  assign T708 = $signed(T710) * $signed(T709);
  assign T709 = 18'h8000;
  assign T710 = T711;
  assign T711 = T1107;
  assign T1107 = T712[5'h11:1'h0];
  assign T712 = $signed(T713) >>> 4'he;
  assign T713 = $signed(T715) * $signed(T714);
  assign T714 = io_lbda;
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = T727 - T718;
  assign T718 = R719;
  assign T727 = R728;
  assign T733 = R734;
  assign io_yout_5 = yout_5;
  assign T737 = T738;
  assign T738 = T770 + T739;
  assign T739 = R740;
  assign T743 = T1108;
  assign T1108 = T744[5'h11:1'h0];
  assign T744 = $signed(T745) >>> 4'he;
  assign T745 = $signed(T747) * $signed(T746);
  assign T746 = 18'h8000;
  assign T747 = T748;
  assign T748 = T1109;
  assign T1109 = T749[5'h11:1'h0];
  assign T749 = $signed(T750) >>> 4'he;
  assign T750 = $signed(T752) * $signed(T751);
  assign T751 = io_lbda;
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T764 - T755;
  assign T755 = R756;
  assign T764 = R765;
  assign T770 = R771;
  assign io_yout_6 = yout_6;
  assign T774 = T775;
  assign T775 = T807 + T776;
  assign T776 = R777;
  assign T780 = T1110;
  assign T1110 = T781[5'h11:1'h0];
  assign T781 = $signed(T782) >>> 4'he;
  assign T782 = $signed(T784) * $signed(T783);
  assign T783 = 18'h8000;
  assign T784 = T785;
  assign T785 = T1111;
  assign T1111 = T786[5'h11:1'h0];
  assign T786 = $signed(T787) >>> 4'he;
  assign T787 = $signed(T789) * $signed(T788);
  assign T788 = io_lbda;
  assign T789 = T790;
  assign T790 = T791;
  assign T791 = T801 - T792;
  assign T792 = R793;
  assign T801 = R802;
  assign T807 = R808;
  assign io_yout_7 = yout_7;
  assign T811 = T812;
  assign T812 = T844 + T813;
  assign T813 = R814;
  assign T817 = T1112;
  assign T1112 = T818[5'h11:1'h0];
  assign T818 = $signed(T819) >>> 4'he;
  assign T819 = $signed(T821) * $signed(T820);
  assign T820 = 18'h8000;
  assign T821 = T822;
  assign T822 = T1113;
  assign T1113 = T823[5'h11:1'h0];
  assign T823 = $signed(T824) >>> 4'he;
  assign T824 = $signed(T826) * $signed(T825);
  assign T825 = io_lbda;
  assign T826 = T827;
  assign T827 = T828;
  assign T828 = T838 - T829;
  assign T829 = R830;
  assign T838 = R839;
  assign T844 = R845;
  assign io_yout_8 = yout_8;
  assign T848 = T849;
  assign T849 = T881 + T850;
  assign T850 = R851;
  assign T854 = T1114;
  assign T1114 = T855[5'h11:1'h0];
  assign T855 = $signed(T856) >>> 4'he;
  assign T856 = $signed(T858) * $signed(T857);
  assign T857 = 18'h8000;
  assign T858 = T859;
  assign T859 = T1115;
  assign T1115 = T860[5'h11:1'h0];
  assign T860 = $signed(T861) >>> 4'he;
  assign T861 = $signed(T863) * $signed(T862);
  assign T862 = io_lbda;
  assign T863 = T864;
  assign T864 = T865;
  assign T865 = T875 - T866;
  assign T866 = R867;
  assign T875 = R876;
  assign T881 = R882;
  assign io_yout_9 = yout_9;
  assign T885 = T886;
  assign T886 = T918 + T887;
  assign T887 = R888;
  assign T891 = T1116;
  assign T1116 = T892[5'h11:1'h0];
  assign T892 = $signed(T893) >>> 4'he;
  assign T893 = $signed(T895) * $signed(T894);
  assign T894 = 18'h8000;
  assign T895 = T896;
  assign T896 = T1117;
  assign T1117 = T897[5'h11:1'h0];
  assign T897 = $signed(T898) >>> 4'he;
  assign T898 = $signed(T900) * $signed(T899);
  assign T899 = io_lbda;
  assign T900 = T901;
  assign T901 = T902;
  assign T902 = T912 - T903;
  assign T903 = R904;
  assign T912 = R913;
  assign T918 = R919;
  assign io_yout_10 = yout_10;
  assign T922 = T923;
  assign T923 = T955 + T924;
  assign T924 = R925;
  assign T928 = T1118;
  assign T1118 = T929[5'h11:1'h0];
  assign T929 = $signed(T930) >>> 4'he;
  assign T930 = $signed(T932) * $signed(T931);
  assign T931 = 18'h8000;
  assign T932 = T933;
  assign T933 = T1119;
  assign T1119 = T934[5'h11:1'h0];
  assign T934 = $signed(T935) >>> 4'he;
  assign T935 = $signed(T937) * $signed(T936);
  assign T936 = io_lbda;
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = T949 - T940;
  assign T940 = R941;
  assign T949 = R950;
  assign T955 = R956;
  assign io_yout_11 = yout_11;
  assign T959 = T960;
  assign T960 = T992 + T961;
  assign T961 = R962;
  assign T965 = T1120;
  assign T1120 = T966[5'h11:1'h0];
  assign T966 = $signed(T967) >>> 4'he;
  assign T967 = $signed(T969) * $signed(T968);
  assign T968 = 18'h8000;
  assign T969 = T970;
  assign T970 = T1121;
  assign T1121 = T971[5'h11:1'h0];
  assign T971 = $signed(T972) >>> 4'he;
  assign T972 = $signed(T974) * $signed(T973);
  assign T973 = io_lbda;
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T986 - T977;
  assign T977 = R978;
  assign T986 = R987;
  assign T992 = R993;
  assign io_xout_0 = xout_0;
  assign T996 = T997;
  assign T997 = T1024 + T998;
  assign T998 = R999;
  assign T1002 = T1122;
  assign T1122 = T1003[5'h11:1'h0];
  assign T1003 = $signed(T1004) >>> 4'he;
  assign T1004 = $signed(T1006) * $signed(T1005);
  assign T1005 = io_lbda;
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1023 - T1009;
  assign T1009 = R1010;
  assign T1023 = R0;
  assign T1024 = R1025;
  assign io_xout_1 = xout_1;
  assign T1028 = T1029;
  assign T1029 = T1056 + T1030;
  assign T1030 = R1031;
  assign T1034 = T1123;
  assign T1123 = T1035[5'h11:1'h0];
  assign T1035 = $signed(T1036) >>> 4'he;
  assign T1036 = $signed(T1038) * $signed(T1037);
  assign T1037 = io_lbda;
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1055 - T1041;
  assign T1041 = R1042;
  assign T1055 = R9;
  assign T1056 = R1057;
  assign io_xout_2 = xout_2;
  assign T1060 = T1061;
  assign T1061 = T1088 + T1062;
  assign T1062 = R1063;
  assign T1066 = T1124;
  assign T1124 = T1067[5'h11:1'h0];
  assign T1067 = $signed(T1068) >>> 4'he;
  assign T1068 = $signed(T1070) * $signed(T1069);
  assign T1069 = io_lbda;
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1087 - T1073;
  assign T1073 = R1074;
  assign T1087 = R18;
  assign T1088 = R1089;
  XNetModule XNetModule(.clk(clk),
       .io_x_2( io_x_2 ),
       .io_x_1( io_x_1 ),
       .io_x_0( io_x_0 ),
       .io_y_11( io_y_11 ),
       .io_y_10( io_y_10 ),
       .io_y_9( io_y_9 ),
       .io_y_8( io_y_8 ),
       .io_y_7( io_y_7 ),
       .io_y_6( io_y_6 ),
       .io_y_5( io_y_5 ),
       .io_y_4( io_y_4 ),
       .io_y_3( io_y_3 ),
       .io_y_2( io_y_2 ),
       .io_y_1( io_y_1 ),
       .io_y_0( io_y_0 ),
       .io_z_2( io_z_2 ),
       .io_z_1( io_z_1 ),
       .io_z_0( io_z_0 ),
       .io_a_11_2( io_a_11_2 ),
       .io_a_11_1( io_a_11_1 ),
       .io_a_11_0( io_a_11_0 ),
       .io_a_10_2( io_a_10_2 ),
       .io_a_10_1( io_a_10_1 ),
       .io_a_10_0( io_a_10_0 ),
       .io_a_9_2( io_a_9_2 ),
       .io_a_9_1( io_a_9_1 ),
       .io_a_9_0( io_a_9_0 ),
       .io_a_8_2( io_a_8_2 ),
       .io_a_8_1( io_a_8_1 ),
       .io_a_8_0( io_a_8_0 ),
       .io_a_7_2( io_a_7_2 ),
       .io_a_7_1( io_a_7_1 ),
       .io_a_7_0( io_a_7_0 ),
       .io_a_6_2( io_a_6_2 ),
       .io_a_6_1( io_a_6_1 ),
       .io_a_6_0( io_a_6_0 ),
       .io_a_5_2( io_a_5_2 ),
       .io_a_5_1( io_a_5_1 ),
       .io_a_5_0( io_a_5_0 ),
       .io_a_4_2( io_a_4_2 ),
       .io_a_4_1( io_a_4_1 ),
       .io_a_4_0( io_a_4_0 ),
       .io_a_3_2( io_a_3_2 ),
       .io_a_3_1( io_a_3_1 ),
       .io_a_3_0( io_a_3_0 ),
       .io_a_2_2( io_a_2_2 ),
       .io_a_2_1( io_a_2_1 ),
       .io_a_2_0( io_a_2_0 ),
       .io_a_1_2( io_a_1_2 ),
       .io_a_1_1( io_a_1_1 ),
       .io_a_1_0( io_a_1_0 ),
       .io_a_0_2( io_a_0_2 ),
       .io_a_0_1( io_a_0_1 ),
       .io_a_0_0( io_a_0_0 ),
       .io_c_2_2( io_c_2_2 ),
       .io_c_2_1( io_c_2_1 ),
       .io_c_2_0( io_c_2_0 ),
       .io_c_1_2( io_c_1_2 ),
       .io_c_1_1( io_c_1_1 ),
       .io_c_1_0( io_c_1_0 ),
       .io_c_0_2( io_c_0_2 ),
       .io_c_0_1( io_c_0_1 ),
       .io_c_0_0( io_c_0_0 ),
       .io_o_2( XNetModule_io_o_2 ),
       .io_o_1( XNetModule_io_o_1 ),
       .io_o_0( XNetModule_io_o_0 )
  );
  YNetModule YNetModule(.clk(clk),
       .io_x_2( R26 ),
       .io_x_1( R17 ),
       .io_x_0( R8 ),
       .io_y_11( R466 ),
       .io_y_10( R461 ),
       .io_y_9( R456 ),
       .io_y_8( R451 ),
       .io_y_7( R446 ),
       .io_y_6( R441 ),
       .io_y_5( R436 ),
       .io_y_4( R431 ),
       .io_y_3( R426 ),
       .io_y_2( R421 ),
       .io_y_1( R416 ),
       .io_y_0( R411 ),
       .io_b_11( R406 ),
       .io_b_10( R401 ),
       .io_b_9( R396 ),
       .io_b_8( R391 ),
       .io_b_7( R386 ),
       .io_b_6( R381 ),
       .io_b_5( R376 ),
       .io_b_4( R371 ),
       .io_b_3( R366 ),
       .io_b_2( R361 ),
       .io_b_1( R356 ),
       .io_b_0( R351 ),
       .io_a_11_2( R346 ),
       .io_a_11_1( R341 ),
       .io_a_11_0( R336 ),
       .io_a_10_2( R331 ),
       .io_a_10_1( R326 ),
       .io_a_10_0( R321 ),
       .io_a_9_2( R316 ),
       .io_a_9_1( R311 ),
       .io_a_9_0( R306 ),
       .io_a_8_2( R301 ),
       .io_a_8_1( R296 ),
       .io_a_8_0( R291 ),
       .io_a_7_2( R286 ),
       .io_a_7_1( R281 ),
       .io_a_7_0( R276 ),
       .io_a_6_2( R271 ),
       .io_a_6_1( R266 ),
       .io_a_6_0( R261 ),
       .io_a_5_2( R256 ),
       .io_a_5_1( R251 ),
       .io_a_5_0( R246 ),
       .io_a_4_2( R241 ),
       .io_a_4_1( R236 ),
       .io_a_4_0( R231 ),
       .io_a_3_2( R226 ),
       .io_a_3_1( R221 ),
       .io_a_3_0( R216 ),
       .io_a_2_2( R211 ),
       .io_a_2_1( R206 ),
       .io_a_2_0( R201 ),
       .io_a_1_2( R196 ),
       .io_a_1_1( R191 ),
       .io_a_1_0( R186 ),
       .io_a_0_2( R181 ),
       .io_a_0_1( R176 ),
       .io_a_0_0( R171 ),
       .io_o_11( YNetModule_io_o_11 ),
       .io_o_10( YNetModule_io_o_10 ),
       .io_o_9( YNetModule_io_o_9 ),
       .io_o_8( YNetModule_io_o_8 ),
       .io_o_7( YNetModule_io_o_7 ),
       .io_o_6( YNetModule_io_o_6 ),
       .io_o_5( YNetModule_io_o_5 ),
       .io_o_4( YNetModule_io_o_4 ),
       .io_o_3( YNetModule_io_o_3 ),
       .io_o_2( YNetModule_io_o_2 ),
       .io_o_1( YNetModule_io_o_1 ),
       .io_o_0( YNetModule_io_o_0 )
  );
  ZNetModule ZNetModule(.clk(clk),
       .io_x_2( R22 ),
       .io_x_1( R13 ),
       .io_x_0( R4 ),
       .io_z_2( R162 ),
       .io_z_1( R153 ),
       .io_z_0( R144 ),
       .io_c_2_2( R135 ),
       .io_c_2_1( R122 ),
       .io_c_2_0( R109 ),
       .io_c_1_2( R96 ),
       .io_c_1_1( R83 ),
       .io_c_1_0( R70 ),
       .io_c_0_2( R57 ),
       .io_c_0_1( R44 ),
       .io_c_0_0( R31 ),
       .io_o_2( ZNetModule_io_o_2 ),
       .io_o_1( ZNetModule_io_o_1 ),
       .io_o_0( ZNetModule_io_o_0 )
  );
  MatrixVectorMultModule_0 MatrixVectorMultModule(.clk(clk),
       .io_a_2_2( R131 ),
       .io_a_2_1( R118 ),
       .io_a_2_0( R105 ),
       .io_a_1_2( R92 ),
       .io_a_1_1( R79 ),
       .io_a_1_0( R66 ),
       .io_a_0_2( R53 ),
       .io_a_0_1( R40 ),
       .io_a_0_0( R27 ),
       .io_b_2( R18 ),
       .io_b_1( R9 ),
       .io_b_0( R0 ),
       .io_o_2( MatrixVectorMultModule_io_o_2 ),
       .io_o_1( MatrixVectorMultModule_io_o_1 ),
       .io_o_0( MatrixVectorMultModule_io_o_0 )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= R2;
    R2 <= R3;
    R3 <= R4;
    R4 <= R5;
    R5 <= R6;
    R6 <= R7;
    R7 <= R8;
    R8 <= XNetModule_io_o_0;
    R9 <= R10;
    R10 <= R11;
    R11 <= R12;
    R12 <= R13;
    R13 <= R14;
    R14 <= R15;
    R15 <= R16;
    R16 <= R17;
    R17 <= XNetModule_io_o_1;
    R18 <= R19;
    R19 <= R20;
    R20 <= R21;
    R21 <= R22;
    R22 <= R23;
    R23 <= R24;
    R24 <= R25;
    R25 <= R26;
    R26 <= XNetModule_io_o_2;
    R27 <= R28;
    R28 <= R29;
    R29 <= R30;
    R30 <= R31;
    R31 <= R32;
    R32 <= R33;
    R33 <= R34;
    R34 <= R35;
    R35 <= R36;
    R36 <= R37;
    R37 <= R38;
    R38 <= R39;
    R39 <= io_c_0_0;
    R40 <= R41;
    R41 <= R42;
    R42 <= R43;
    R43 <= R44;
    R44 <= R45;
    R45 <= R46;
    R46 <= R47;
    R47 <= R48;
    R48 <= R49;
    R49 <= R50;
    R50 <= R51;
    R51 <= R52;
    R52 <= io_c_0_1;
    R53 <= R54;
    R54 <= R55;
    R55 <= R56;
    R56 <= R57;
    R57 <= R58;
    R58 <= R59;
    R59 <= R60;
    R60 <= R61;
    R61 <= R62;
    R62 <= R63;
    R63 <= R64;
    R64 <= R65;
    R65 <= io_c_0_2;
    R66 <= R67;
    R67 <= R68;
    R68 <= R69;
    R69 <= R70;
    R70 <= R71;
    R71 <= R72;
    R72 <= R73;
    R73 <= R74;
    R74 <= R75;
    R75 <= R76;
    R76 <= R77;
    R77 <= R78;
    R78 <= io_c_1_0;
    R79 <= R80;
    R80 <= R81;
    R81 <= R82;
    R82 <= R83;
    R83 <= R84;
    R84 <= R85;
    R85 <= R86;
    R86 <= R87;
    R87 <= R88;
    R88 <= R89;
    R89 <= R90;
    R90 <= R91;
    R91 <= io_c_1_1;
    R92 <= R93;
    R93 <= R94;
    R94 <= R95;
    R95 <= R96;
    R96 <= R97;
    R97 <= R98;
    R98 <= R99;
    R99 <= R100;
    R100 <= R101;
    R101 <= R102;
    R102 <= R103;
    R103 <= R104;
    R104 <= io_c_1_2;
    R105 <= R106;
    R106 <= R107;
    R107 <= R108;
    R108 <= R109;
    R109 <= R110;
    R110 <= R111;
    R111 <= R112;
    R112 <= R113;
    R113 <= R114;
    R114 <= R115;
    R115 <= R116;
    R116 <= R117;
    R117 <= io_c_2_0;
    R118 <= R119;
    R119 <= R120;
    R120 <= R121;
    R121 <= R122;
    R122 <= R123;
    R123 <= R124;
    R124 <= R125;
    R125 <= R126;
    R126 <= R127;
    R127 <= R128;
    R128 <= R129;
    R129 <= R130;
    R130 <= io_c_2_1;
    R131 <= R132;
    R132 <= R133;
    R133 <= R134;
    R134 <= R135;
    R135 <= R136;
    R136 <= R137;
    R137 <= R138;
    R138 <= R139;
    R139 <= R140;
    R140 <= R141;
    R141 <= R142;
    R142 <= R143;
    R143 <= io_c_2_2;
    R144 <= R145;
    R145 <= R146;
    R146 <= R147;
    R147 <= R148;
    R148 <= R149;
    R149 <= R150;
    R150 <= R151;
    R151 <= R152;
    R152 <= io_z_0;
    R153 <= R154;
    R154 <= R155;
    R155 <= R156;
    R156 <= R157;
    R157 <= R158;
    R158 <= R159;
    R159 <= R160;
    R160 <= R161;
    R161 <= io_z_1;
    R162 <= R163;
    R163 <= R164;
    R164 <= R165;
    R165 <= R166;
    R166 <= R167;
    R167 <= R168;
    R168 <= R169;
    R169 <= R170;
    R170 <= io_z_2;
    R171 <= R172;
    R172 <= R173;
    R173 <= R174;
    R174 <= R175;
    R175 <= io_a_0_0;
    R176 <= R177;
    R177 <= R178;
    R178 <= R179;
    R179 <= R180;
    R180 <= io_a_0_1;
    R181 <= R182;
    R182 <= R183;
    R183 <= R184;
    R184 <= R185;
    R185 <= io_a_0_2;
    R186 <= R187;
    R187 <= R188;
    R188 <= R189;
    R189 <= R190;
    R190 <= io_a_1_0;
    R191 <= R192;
    R192 <= R193;
    R193 <= R194;
    R194 <= R195;
    R195 <= io_a_1_1;
    R196 <= R197;
    R197 <= R198;
    R198 <= R199;
    R199 <= R200;
    R200 <= io_a_1_2;
    R201 <= R202;
    R202 <= R203;
    R203 <= R204;
    R204 <= R205;
    R205 <= io_a_2_0;
    R206 <= R207;
    R207 <= R208;
    R208 <= R209;
    R209 <= R210;
    R210 <= io_a_2_1;
    R211 <= R212;
    R212 <= R213;
    R213 <= R214;
    R214 <= R215;
    R215 <= io_a_2_2;
    R216 <= R217;
    R217 <= R218;
    R218 <= R219;
    R219 <= R220;
    R220 <= io_a_3_0;
    R221 <= R222;
    R222 <= R223;
    R223 <= R224;
    R224 <= R225;
    R225 <= io_a_3_1;
    R226 <= R227;
    R227 <= R228;
    R228 <= R229;
    R229 <= R230;
    R230 <= io_a_3_2;
    R231 <= R232;
    R232 <= R233;
    R233 <= R234;
    R234 <= R235;
    R235 <= io_a_4_0;
    R236 <= R237;
    R237 <= R238;
    R238 <= R239;
    R239 <= R240;
    R240 <= io_a_4_1;
    R241 <= R242;
    R242 <= R243;
    R243 <= R244;
    R244 <= R245;
    R245 <= io_a_4_2;
    R246 <= R247;
    R247 <= R248;
    R248 <= R249;
    R249 <= R250;
    R250 <= io_a_5_0;
    R251 <= R252;
    R252 <= R253;
    R253 <= R254;
    R254 <= R255;
    R255 <= io_a_5_1;
    R256 <= R257;
    R257 <= R258;
    R258 <= R259;
    R259 <= R260;
    R260 <= io_a_5_2;
    R261 <= R262;
    R262 <= R263;
    R263 <= R264;
    R264 <= R265;
    R265 <= io_a_6_0;
    R266 <= R267;
    R267 <= R268;
    R268 <= R269;
    R269 <= R270;
    R270 <= io_a_6_1;
    R271 <= R272;
    R272 <= R273;
    R273 <= R274;
    R274 <= R275;
    R275 <= io_a_6_2;
    R276 <= R277;
    R277 <= R278;
    R278 <= R279;
    R279 <= R280;
    R280 <= io_a_7_0;
    R281 <= R282;
    R282 <= R283;
    R283 <= R284;
    R284 <= R285;
    R285 <= io_a_7_1;
    R286 <= R287;
    R287 <= R288;
    R288 <= R289;
    R289 <= R290;
    R290 <= io_a_7_2;
    R291 <= R292;
    R292 <= R293;
    R293 <= R294;
    R294 <= R295;
    R295 <= io_a_8_0;
    R296 <= R297;
    R297 <= R298;
    R298 <= R299;
    R299 <= R300;
    R300 <= io_a_8_1;
    R301 <= R302;
    R302 <= R303;
    R303 <= R304;
    R304 <= R305;
    R305 <= io_a_8_2;
    R306 <= R307;
    R307 <= R308;
    R308 <= R309;
    R309 <= R310;
    R310 <= io_a_9_0;
    R311 <= R312;
    R312 <= R313;
    R313 <= R314;
    R314 <= R315;
    R315 <= io_a_9_1;
    R316 <= R317;
    R317 <= R318;
    R318 <= R319;
    R319 <= R320;
    R320 <= io_a_9_2;
    R321 <= R322;
    R322 <= R323;
    R323 <= R324;
    R324 <= R325;
    R325 <= io_a_10_0;
    R326 <= R327;
    R327 <= R328;
    R328 <= R329;
    R329 <= R330;
    R330 <= io_a_10_1;
    R331 <= R332;
    R332 <= R333;
    R333 <= R334;
    R334 <= R335;
    R335 <= io_a_10_2;
    R336 <= R337;
    R337 <= R338;
    R338 <= R339;
    R339 <= R340;
    R340 <= io_a_11_0;
    R341 <= R342;
    R342 <= R343;
    R343 <= R344;
    R344 <= R345;
    R345 <= io_a_11_1;
    R346 <= R347;
    R347 <= R348;
    R348 <= R349;
    R349 <= R350;
    R350 <= io_a_11_2;
    R351 <= R352;
    R352 <= R353;
    R353 <= R354;
    R354 <= R355;
    R355 <= io_b_0;
    R356 <= R357;
    R357 <= R358;
    R358 <= R359;
    R359 <= R360;
    R360 <= io_b_1;
    R361 <= R362;
    R362 <= R363;
    R363 <= R364;
    R364 <= R365;
    R365 <= io_b_2;
    R366 <= R367;
    R367 <= R368;
    R368 <= R369;
    R369 <= R370;
    R370 <= io_b_3;
    R371 <= R372;
    R372 <= R373;
    R373 <= R374;
    R374 <= R375;
    R375 <= io_b_4;
    R376 <= R377;
    R377 <= R378;
    R378 <= R379;
    R379 <= R380;
    R380 <= io_b_5;
    R381 <= R382;
    R382 <= R383;
    R383 <= R384;
    R384 <= R385;
    R385 <= io_b_6;
    R386 <= R387;
    R387 <= R388;
    R388 <= R389;
    R389 <= R390;
    R390 <= io_b_7;
    R391 <= R392;
    R392 <= R393;
    R393 <= R394;
    R394 <= R395;
    R395 <= io_b_8;
    R396 <= R397;
    R397 <= R398;
    R398 <= R399;
    R399 <= R400;
    R400 <= io_b_9;
    R401 <= R402;
    R402 <= R403;
    R403 <= R404;
    R404 <= R405;
    R405 <= io_b_10;
    R406 <= R407;
    R407 <= R408;
    R408 <= R409;
    R409 <= R410;
    R410 <= io_b_11;
    R411 <= R412;
    R412 <= R413;
    R413 <= R414;
    R414 <= R415;
    R415 <= io_y_0;
    R416 <= R417;
    R417 <= R418;
    R418 <= R419;
    R419 <= R420;
    R420 <= io_y_1;
    R421 <= R422;
    R422 <= R423;
    R423 <= R424;
    R424 <= R425;
    R425 <= io_y_2;
    R426 <= R427;
    R427 <= R428;
    R428 <= R429;
    R429 <= R430;
    R430 <= io_y_3;
    R431 <= R432;
    R432 <= R433;
    R433 <= R434;
    R434 <= R435;
    R435 <= io_y_4;
    R436 <= R437;
    R437 <= R438;
    R438 <= R439;
    R439 <= R440;
    R440 <= io_y_5;
    R441 <= R442;
    R442 <= R443;
    R443 <= R444;
    R444 <= R445;
    R445 <= io_y_6;
    R446 <= R447;
    R447 <= R448;
    R448 <= R449;
    R449 <= R450;
    R450 <= io_y_7;
    R451 <= R452;
    R452 <= R453;
    R453 <= R454;
    R454 <= R455;
    R455 <= io_y_8;
    R456 <= R457;
    R457 <= R458;
    R458 <= R459;
    R459 <= R460;
    R460 <= io_y_9;
    R461 <= R462;
    R462 <= R463;
    R463 <= R464;
    R464 <= R465;
    R465 <= io_y_10;
    R466 <= R467;
    R467 <= R468;
    R468 <= R469;
    R469 <= R470;
    R470 <= io_y_11;
    zout_0 <= T471;
    R474 <= T475;
    R488 <= ZNetModule_io_o_0;
    R491 <= R492;
    R492 <= R493;
    R493 <= R494;
    R494 <= R495;
    R495 <= R496;
    R496 <= R497;
    R497 <= R144;
    zout_1 <= T498;
    R501 <= T502;
    R515 <= ZNetModule_io_o_1;
    R518 <= R519;
    R519 <= R520;
    R520 <= R521;
    R521 <= R522;
    R522 <= R523;
    R523 <= R524;
    R524 <= R153;
    zout_2 <= T525;
    R528 <= T529;
    R542 <= ZNetModule_io_o_2;
    R545 <= R546;
    R546 <= R547;
    R547 <= R548;
    R548 <= R549;
    R549 <= R550;
    R550 <= R551;
    R551 <= R162;
    yout_0 <= T552;
    R555 <= R556;
    R556 <= R557;
    R557 <= T558;
    R571 <= R572;
    R572 <= R573;
    R573 <= R574;
    R574 <= R575;
    R575 <= R576;
    R576 <= R577;
    R577 <= R578;
    R578 <= R411;
    R580 <= R581;
    R581 <= R582;
    R582 <= R583;
    R583 <= R584;
    R584 <= YNetModule_io_o_0;
    R586 <= R587;
    R587 <= R588;
    R588 <= R571;
    yout_1 <= T589;
    R592 <= R593;
    R593 <= R594;
    R594 <= T595;
    R608 <= R609;
    R609 <= R610;
    R610 <= R611;
    R611 <= R612;
    R612 <= R613;
    R613 <= R614;
    R614 <= R615;
    R615 <= R416;
    R617 <= R618;
    R618 <= R619;
    R619 <= R620;
    R620 <= R621;
    R621 <= YNetModule_io_o_1;
    R623 <= R624;
    R624 <= R625;
    R625 <= R608;
    yout_2 <= T626;
    R629 <= R630;
    R630 <= R631;
    R631 <= T632;
    R645 <= R646;
    R646 <= R647;
    R647 <= R648;
    R648 <= R649;
    R649 <= R650;
    R650 <= R651;
    R651 <= R652;
    R652 <= R421;
    R654 <= R655;
    R655 <= R656;
    R656 <= R657;
    R657 <= R658;
    R658 <= YNetModule_io_o_2;
    R660 <= R661;
    R661 <= R662;
    R662 <= R645;
    yout_3 <= T663;
    R666 <= R667;
    R667 <= R668;
    R668 <= T669;
    R682 <= R683;
    R683 <= R684;
    R684 <= R685;
    R685 <= R686;
    R686 <= R687;
    R687 <= R688;
    R688 <= R689;
    R689 <= R426;
    R691 <= R692;
    R692 <= R693;
    R693 <= R694;
    R694 <= R695;
    R695 <= YNetModule_io_o_3;
    R697 <= R698;
    R698 <= R699;
    R699 <= R682;
    yout_4 <= T700;
    R703 <= R704;
    R704 <= R705;
    R705 <= T706;
    R719 <= R720;
    R720 <= R721;
    R721 <= R722;
    R722 <= R723;
    R723 <= R724;
    R724 <= R725;
    R725 <= R726;
    R726 <= R431;
    R728 <= R729;
    R729 <= R730;
    R730 <= R731;
    R731 <= R732;
    R732 <= YNetModule_io_o_4;
    R734 <= R735;
    R735 <= R736;
    R736 <= R719;
    yout_5 <= T737;
    R740 <= R741;
    R741 <= R742;
    R742 <= T743;
    R756 <= R757;
    R757 <= R758;
    R758 <= R759;
    R759 <= R760;
    R760 <= R761;
    R761 <= R762;
    R762 <= R763;
    R763 <= R436;
    R765 <= R766;
    R766 <= R767;
    R767 <= R768;
    R768 <= R769;
    R769 <= YNetModule_io_o_5;
    R771 <= R772;
    R772 <= R773;
    R773 <= R756;
    yout_6 <= T774;
    R777 <= R778;
    R778 <= R779;
    R779 <= T780;
    R793 <= R794;
    R794 <= R795;
    R795 <= R796;
    R796 <= R797;
    R797 <= R798;
    R798 <= R799;
    R799 <= R800;
    R800 <= R441;
    R802 <= R803;
    R803 <= R804;
    R804 <= R805;
    R805 <= R806;
    R806 <= YNetModule_io_o_6;
    R808 <= R809;
    R809 <= R810;
    R810 <= R793;
    yout_7 <= T811;
    R814 <= R815;
    R815 <= R816;
    R816 <= T817;
    R830 <= R831;
    R831 <= R832;
    R832 <= R833;
    R833 <= R834;
    R834 <= R835;
    R835 <= R836;
    R836 <= R837;
    R837 <= R446;
    R839 <= R840;
    R840 <= R841;
    R841 <= R842;
    R842 <= R843;
    R843 <= YNetModule_io_o_7;
    R845 <= R846;
    R846 <= R847;
    R847 <= R830;
    yout_8 <= T848;
    R851 <= R852;
    R852 <= R853;
    R853 <= T854;
    R867 <= R868;
    R868 <= R869;
    R869 <= R870;
    R870 <= R871;
    R871 <= R872;
    R872 <= R873;
    R873 <= R874;
    R874 <= R451;
    R876 <= R877;
    R877 <= R878;
    R878 <= R879;
    R879 <= R880;
    R880 <= YNetModule_io_o_8;
    R882 <= R883;
    R883 <= R884;
    R884 <= R867;
    yout_9 <= T885;
    R888 <= R889;
    R889 <= R890;
    R890 <= T891;
    R904 <= R905;
    R905 <= R906;
    R906 <= R907;
    R907 <= R908;
    R908 <= R909;
    R909 <= R910;
    R910 <= R911;
    R911 <= R456;
    R913 <= R914;
    R914 <= R915;
    R915 <= R916;
    R916 <= R917;
    R917 <= YNetModule_io_o_9;
    R919 <= R920;
    R920 <= R921;
    R921 <= R904;
    yout_10 <= T922;
    R925 <= R926;
    R926 <= R927;
    R927 <= T928;
    R941 <= R942;
    R942 <= R943;
    R943 <= R944;
    R944 <= R945;
    R945 <= R946;
    R946 <= R947;
    R947 <= R948;
    R948 <= R461;
    R950 <= R951;
    R951 <= R952;
    R952 <= R953;
    R953 <= R954;
    R954 <= YNetModule_io_o_10;
    R956 <= R957;
    R957 <= R958;
    R958 <= R941;
    yout_11 <= T959;
    R962 <= R963;
    R963 <= R964;
    R964 <= T965;
    R978 <= R979;
    R979 <= R980;
    R980 <= R981;
    R981 <= R982;
    R982 <= R983;
    R983 <= R984;
    R984 <= R985;
    R985 <= R466;
    R987 <= R988;
    R988 <= R989;
    R989 <= R990;
    R990 <= R991;
    R991 <= YNetModule_io_o_11;
    R993 <= R994;
    R994 <= R995;
    R995 <= R978;
    xout_0 <= T996;
    R999 <= R1000;
    R1000 <= R1001;
    R1001 <= T1002;
    R1010 <= R1011;
    R1011 <= R1012;
    R1012 <= R1013;
    R1013 <= R1014;
    R1014 <= R1015;
    R1015 <= R1016;
    R1016 <= R1017;
    R1017 <= R1018;
    R1018 <= R1019;
    R1019 <= R1020;
    R1020 <= R1021;
    R1021 <= R1022;
    R1022 <= io_x_0;
    R1025 <= R1026;
    R1026 <= R1027;
    R1027 <= R1010;
    xout_1 <= T1028;
    R1031 <= R1032;
    R1032 <= R1033;
    R1033 <= T1034;
    R1042 <= R1043;
    R1043 <= R1044;
    R1044 <= R1045;
    R1045 <= R1046;
    R1046 <= R1047;
    R1047 <= R1048;
    R1048 <= R1049;
    R1049 <= R1050;
    R1050 <= R1051;
    R1051 <= R1052;
    R1052 <= R1053;
    R1053 <= R1054;
    R1054 <= io_x_1;
    R1057 <= R1058;
    R1058 <= R1059;
    R1059 <= R1042;
    xout_2 <= T1060;
    R1063 <= R1064;
    R1064 <= R1065;
    R1065 <= T1066;
    R1074 <= R1075;
    R1075 <= R1076;
    R1076 <= R1077;
    R1077 <= R1078;
    R1078 <= R1079;
    R1079 <= R1080;
    R1080 <= R1081;
    R1081 <= R1082;
    R1082 <= R1083;
    R1083 <= R1084;
    R1084 <= R1085;
    R1085 <= R1086;
    R1086 <= io_x_2;
    R1089 <= R1090;
    R1090 <= R1091;
    R1091 <= R1074;
  end
endmodule

module NN1ShiftTop(input clk, input reset,
    input [17:0] io_x,
    input [17:0] io_y,
    input [17:0] io_z,
    input [17:0] io_b,
    input [17:0] io_a,
    input [17:0] io_c,
    input [17:0] io_lbda,
    output[17:0] io_xout,
    output[17:0] io_yout,
    output[17:0] io_zout
);

  reg [17:0] cShift_0_0;
  wire[17:0] T60;
  reg [17:0] cShift_1_0;
  wire[17:0] T61;
  reg [17:0] cShift_2_0;
  wire[17:0] T62;
  reg [17:0] cShift_0_1;
  wire[17:0] T63;
  reg [17:0] cShift_1_1;
  wire[17:0] T64;
  reg [17:0] cShift_2_1;
  wire[17:0] T65;
  reg [17:0] cShift_0_2;
  wire[17:0] T66;
  reg [17:0] cShift_1_2;
  wire[17:0] T67;
  reg [17:0] cShift_2_2;
  wire[17:0] T68;
  reg [17:0] aShift_0_0;
  wire[17:0] T69;
  reg [17:0] aShift_1_0;
  wire[17:0] T70;
  reg [17:0] aShift_2_0;
  wire[17:0] T71;
  reg [17:0] aShift_3_0;
  wire[17:0] T72;
  reg [17:0] aShift_4_0;
  wire[17:0] T73;
  reg [17:0] aShift_5_0;
  wire[17:0] T74;
  reg [17:0] aShift_6_0;
  wire[17:0] T75;
  reg [17:0] aShift_7_0;
  wire[17:0] T76;
  reg [17:0] aShift_8_0;
  wire[17:0] T77;
  reg [17:0] aShift_9_0;
  wire[17:0] T78;
  reg [17:0] aShift_10_0;
  wire[17:0] T79;
  reg [17:0] aShift_11_0;
  wire[17:0] T80;
  reg [17:0] aShift_0_1;
  wire[17:0] T81;
  reg [17:0] aShift_1_1;
  wire[17:0] T82;
  reg [17:0] aShift_2_1;
  wire[17:0] T83;
  reg [17:0] aShift_3_1;
  wire[17:0] T84;
  reg [17:0] aShift_4_1;
  wire[17:0] T85;
  reg [17:0] aShift_5_1;
  wire[17:0] T86;
  reg [17:0] aShift_6_1;
  wire[17:0] T87;
  reg [17:0] aShift_7_1;
  wire[17:0] T88;
  reg [17:0] aShift_8_1;
  wire[17:0] T89;
  reg [17:0] aShift_9_1;
  wire[17:0] T90;
  reg [17:0] aShift_10_1;
  wire[17:0] T91;
  reg [17:0] aShift_11_1;
  wire[17:0] T92;
  reg [17:0] aShift_0_2;
  wire[17:0] T93;
  reg [17:0] aShift_1_2;
  wire[17:0] T94;
  reg [17:0] aShift_2_2;
  wire[17:0] T95;
  reg [17:0] aShift_3_2;
  wire[17:0] T96;
  reg [17:0] aShift_4_2;
  wire[17:0] T97;
  reg [17:0] aShift_5_2;
  wire[17:0] T98;
  reg [17:0] aShift_6_2;
  wire[17:0] T99;
  reg [17:0] aShift_7_2;
  wire[17:0] T100;
  reg [17:0] aShift_8_2;
  wire[17:0] T101;
  reg [17:0] aShift_9_2;
  wire[17:0] T102;
  reg [17:0] aShift_10_2;
  wire[17:0] T103;
  reg [17:0] aShift_11_2;
  wire[17:0] T104;
  reg [17:0] bShift_0;
  wire[17:0] T105;
  reg [17:0] bShift_1;
  wire[17:0] T106;
  reg [17:0] bShift_2;
  wire[17:0] T107;
  reg [17:0] bShift_3;
  wire[17:0] T108;
  reg [17:0] bShift_4;
  wire[17:0] T109;
  reg [17:0] bShift_5;
  wire[17:0] T110;
  reg [17:0] bShift_6;
  wire[17:0] T111;
  reg [17:0] bShift_7;
  wire[17:0] T112;
  reg [17:0] bShift_8;
  wire[17:0] T113;
  reg [17:0] bShift_9;
  wire[17:0] T114;
  reg [17:0] bShift_10;
  wire[17:0] T115;
  reg [17:0] bShift_11;
  wire[17:0] T116;
  reg [17:0] zShift_0;
  wire[17:0] T117;
  reg [17:0] zShift_1;
  wire[17:0] T118;
  reg [17:0] zShift_2;
  wire[17:0] T119;
  reg [17:0] yShift_0;
  wire[17:0] T120;
  reg [17:0] yShift_1;
  wire[17:0] T121;
  reg [17:0] yShift_2;
  wire[17:0] T122;
  reg [17:0] yShift_3;
  wire[17:0] T123;
  reg [17:0] yShift_4;
  wire[17:0] T124;
  reg [17:0] yShift_5;
  wire[17:0] T125;
  reg [17:0] yShift_6;
  wire[17:0] T126;
  reg [17:0] yShift_7;
  wire[17:0] T127;
  reg [17:0] yShift_8;
  wire[17:0] T128;
  reg [17:0] yShift_9;
  wire[17:0] T129;
  reg [17:0] yShift_10;
  wire[17:0] T130;
  reg [17:0] yShift_11;
  wire[17:0] T131;
  reg [17:0] xShift_0;
  wire[17:0] T132;
  reg [17:0] xShift_1;
  wire[17:0] T133;
  reg [17:0] xShift_2;
  wire[17:0] T134;
  reg [17:0] nnzout;
  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  wire[17:0] T3;
  wire[17:0] T4;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  reg [17:0] nnyout;
  wire[17:0] T8;
  wire[17:0] T9;
  wire[17:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  wire[17:0] T16;
  wire[17:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  wire[17:0] T20;
  wire[17:0] T21;
  wire[17:0] T22;
  wire[17:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;
  wire[17:0] T26;
  wire[17:0] T27;
  wire[17:0] T28;
  wire[17:0] T29;
  wire[17:0] T30;
  wire[17:0] T31;
  wire[17:0] T32;
  wire[17:0] T33;
  wire[17:0] T34;
  wire[17:0] T35;
  wire[17:0] T36;
  wire[17:0] T37;
  wire[17:0] T38;
  wire[17:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  wire[17:0] T42;
  wire[17:0] T43;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[17:0] T46;
  wire[17:0] T47;
  wire[17:0] T48;
  wire[17:0] T49;
  wire[17:0] T50;
  wire[17:0] T51;
  reg [17:0] nnxout;
  wire[17:0] T52;
  wire[17:0] T53;
  wire[17:0] T54;
  wire[17:0] T55;
  wire[17:0] T56;
  wire[17:0] T57;
  wire[17:0] T58;
  wire[17:0] T59;
  wire[17:0] nnTop_io_xout_2;
  wire[17:0] nnTop_io_xout_1;
  wire[17:0] nnTop_io_xout_0;
  wire[17:0] nnTop_io_yout_11;
  wire[17:0] nnTop_io_yout_10;
  wire[17:0] nnTop_io_yout_9;
  wire[17:0] nnTop_io_yout_8;
  wire[17:0] nnTop_io_yout_7;
  wire[17:0] nnTop_io_yout_6;
  wire[17:0] nnTop_io_yout_5;
  wire[17:0] nnTop_io_yout_4;
  wire[17:0] nnTop_io_yout_3;
  wire[17:0] nnTop_io_yout_2;
  wire[17:0] nnTop_io_yout_1;
  wire[17:0] nnTop_io_yout_0;
  wire[17:0] nnTop_io_zout_2;
  wire[17:0] nnTop_io_zout_1;
  wire[17:0] nnTop_io_zout_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    cShift_0_0 = {1{$random}};
    cShift_1_0 = {1{$random}};
    cShift_2_0 = {1{$random}};
    cShift_0_1 = {1{$random}};
    cShift_1_1 = {1{$random}};
    cShift_2_1 = {1{$random}};
    cShift_0_2 = {1{$random}};
    cShift_1_2 = {1{$random}};
    cShift_2_2 = {1{$random}};
    aShift_0_0 = {1{$random}};
    aShift_1_0 = {1{$random}};
    aShift_2_0 = {1{$random}};
    aShift_3_0 = {1{$random}};
    aShift_4_0 = {1{$random}};
    aShift_5_0 = {1{$random}};
    aShift_6_0 = {1{$random}};
    aShift_7_0 = {1{$random}};
    aShift_8_0 = {1{$random}};
    aShift_9_0 = {1{$random}};
    aShift_10_0 = {1{$random}};
    aShift_11_0 = {1{$random}};
    aShift_0_1 = {1{$random}};
    aShift_1_1 = {1{$random}};
    aShift_2_1 = {1{$random}};
    aShift_3_1 = {1{$random}};
    aShift_4_1 = {1{$random}};
    aShift_5_1 = {1{$random}};
    aShift_6_1 = {1{$random}};
    aShift_7_1 = {1{$random}};
    aShift_8_1 = {1{$random}};
    aShift_9_1 = {1{$random}};
    aShift_10_1 = {1{$random}};
    aShift_11_1 = {1{$random}};
    aShift_0_2 = {1{$random}};
    aShift_1_2 = {1{$random}};
    aShift_2_2 = {1{$random}};
    aShift_3_2 = {1{$random}};
    aShift_4_2 = {1{$random}};
    aShift_5_2 = {1{$random}};
    aShift_6_2 = {1{$random}};
    aShift_7_2 = {1{$random}};
    aShift_8_2 = {1{$random}};
    aShift_9_2 = {1{$random}};
    aShift_10_2 = {1{$random}};
    aShift_11_2 = {1{$random}};
    bShift_0 = {1{$random}};
    bShift_1 = {1{$random}};
    bShift_2 = {1{$random}};
    bShift_3 = {1{$random}};
    bShift_4 = {1{$random}};
    bShift_5 = {1{$random}};
    bShift_6 = {1{$random}};
    bShift_7 = {1{$random}};
    bShift_8 = {1{$random}};
    bShift_9 = {1{$random}};
    bShift_10 = {1{$random}};
    bShift_11 = {1{$random}};
    zShift_0 = {1{$random}};
    zShift_1 = {1{$random}};
    zShift_2 = {1{$random}};
    yShift_0 = {1{$random}};
    yShift_1 = {1{$random}};
    yShift_2 = {1{$random}};
    yShift_3 = {1{$random}};
    yShift_4 = {1{$random}};
    yShift_5 = {1{$random}};
    yShift_6 = {1{$random}};
    yShift_7 = {1{$random}};
    yShift_8 = {1{$random}};
    yShift_9 = {1{$random}};
    yShift_10 = {1{$random}};
    yShift_11 = {1{$random}};
    xShift_0 = {1{$random}};
    xShift_1 = {1{$random}};
    xShift_2 = {1{$random}};
    nnzout = {1{$random}};
    nnyout = {1{$random}};
    nnxout = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T60 = reset ? 18'h0 : cShift_1_0;
  assign T61 = reset ? 18'h0 : cShift_2_0;
  assign T62 = reset ? 18'h0 : io_c;
  assign T63 = reset ? 18'h0 : cShift_1_1;
  assign T64 = reset ? 18'h0 : cShift_2_1;
  assign T65 = reset ? 18'h0 : io_c;
  assign T66 = reset ? 18'h0 : cShift_1_2;
  assign T67 = reset ? 18'h0 : cShift_2_2;
  assign T68 = reset ? 18'h0 : io_c;
  assign T69 = reset ? 18'h0 : aShift_1_0;
  assign T70 = reset ? 18'h0 : aShift_2_0;
  assign T71 = reset ? 18'h0 : aShift_3_0;
  assign T72 = reset ? 18'h0 : aShift_4_0;
  assign T73 = reset ? 18'h0 : aShift_5_0;
  assign T74 = reset ? 18'h0 : aShift_6_0;
  assign T75 = reset ? 18'h0 : aShift_7_0;
  assign T76 = reset ? 18'h0 : aShift_8_0;
  assign T77 = reset ? 18'h0 : aShift_9_0;
  assign T78 = reset ? 18'h0 : aShift_10_0;
  assign T79 = reset ? 18'h0 : aShift_11_0;
  assign T80 = reset ? 18'h0 : io_a;
  assign T81 = reset ? 18'h0 : aShift_1_1;
  assign T82 = reset ? 18'h0 : aShift_2_1;
  assign T83 = reset ? 18'h0 : aShift_3_1;
  assign T84 = reset ? 18'h0 : aShift_4_1;
  assign T85 = reset ? 18'h0 : aShift_5_1;
  assign T86 = reset ? 18'h0 : aShift_6_1;
  assign T87 = reset ? 18'h0 : aShift_7_1;
  assign T88 = reset ? 18'h0 : aShift_8_1;
  assign T89 = reset ? 18'h0 : aShift_9_1;
  assign T90 = reset ? 18'h0 : aShift_10_1;
  assign T91 = reset ? 18'h0 : aShift_11_1;
  assign T92 = reset ? 18'h0 : io_a;
  assign T93 = reset ? 18'h0 : aShift_1_2;
  assign T94 = reset ? 18'h0 : aShift_2_2;
  assign T95 = reset ? 18'h0 : aShift_3_2;
  assign T96 = reset ? 18'h0 : aShift_4_2;
  assign T97 = reset ? 18'h0 : aShift_5_2;
  assign T98 = reset ? 18'h0 : aShift_6_2;
  assign T99 = reset ? 18'h0 : aShift_7_2;
  assign T100 = reset ? 18'h0 : aShift_8_2;
  assign T101 = reset ? 18'h0 : aShift_9_2;
  assign T102 = reset ? 18'h0 : aShift_10_2;
  assign T103 = reset ? 18'h0 : aShift_11_2;
  assign T104 = reset ? 18'h0 : io_a;
  assign T105 = reset ? 18'h0 : bShift_1;
  assign T106 = reset ? 18'h0 : bShift_2;
  assign T107 = reset ? 18'h0 : bShift_3;
  assign T108 = reset ? 18'h0 : bShift_4;
  assign T109 = reset ? 18'h0 : bShift_5;
  assign T110 = reset ? 18'h0 : bShift_6;
  assign T111 = reset ? 18'h0 : bShift_7;
  assign T112 = reset ? 18'h0 : bShift_8;
  assign T113 = reset ? 18'h0 : bShift_9;
  assign T114 = reset ? 18'h0 : bShift_10;
  assign T115 = reset ? 18'h0 : bShift_11;
  assign T116 = reset ? 18'h0 : io_b;
  assign T117 = reset ? 18'h0 : zShift_1;
  assign T118 = reset ? 18'h0 : zShift_2;
  assign T119 = reset ? 18'h0 : io_z;
  assign T120 = reset ? 18'h0 : yShift_1;
  assign T121 = reset ? 18'h0 : yShift_2;
  assign T122 = reset ? 18'h0 : yShift_3;
  assign T123 = reset ? 18'h0 : yShift_4;
  assign T124 = reset ? 18'h0 : yShift_5;
  assign T125 = reset ? 18'h0 : yShift_6;
  assign T126 = reset ? 18'h0 : yShift_7;
  assign T127 = reset ? 18'h0 : yShift_8;
  assign T128 = reset ? 18'h0 : yShift_9;
  assign T129 = reset ? 18'h0 : yShift_10;
  assign T130 = reset ? 18'h0 : yShift_11;
  assign T131 = reset ? 18'h0 : io_y;
  assign T132 = reset ? 18'h0 : xShift_1;
  assign T133 = reset ? 18'h0 : xShift_2;
  assign T134 = reset ? 18'h0 : io_x;
  assign io_zout = nnzout;
  assign T0 = T1;
  assign T1 = T3 + T2;
  assign T2 = nnTop_io_zout_2;
  assign T3 = T4;
  assign T4 = T5;
  assign T5 = T7 + T6;
  assign T6 = nnTop_io_zout_1;
  assign T7 = nnTop_io_zout_0;
  assign io_yout = nnyout;
  assign T8 = T9;
  assign T9 = T11 + T10;
  assign T10 = nnTop_io_yout_11;
  assign T11 = T12;
  assign T12 = T13;
  assign T13 = T15 + T14;
  assign T14 = nnTop_io_yout_10;
  assign T15 = T16;
  assign T16 = T17;
  assign T17 = T19 + T18;
  assign T18 = nnTop_io_yout_9;
  assign T19 = T20;
  assign T20 = T21;
  assign T21 = T23 + T22;
  assign T22 = nnTop_io_yout_8;
  assign T23 = T24;
  assign T24 = T25;
  assign T25 = T27 + T26;
  assign T26 = nnTop_io_yout_7;
  assign T27 = T28;
  assign T28 = T29;
  assign T29 = T31 + T30;
  assign T30 = nnTop_io_yout_6;
  assign T31 = T32;
  assign T32 = T33;
  assign T33 = T35 + T34;
  assign T34 = nnTop_io_yout_5;
  assign T35 = T36;
  assign T36 = T37;
  assign T37 = T39 + T38;
  assign T38 = nnTop_io_yout_4;
  assign T39 = T40;
  assign T40 = T41;
  assign T41 = T43 + T42;
  assign T42 = nnTop_io_yout_3;
  assign T43 = T44;
  assign T44 = T45;
  assign T45 = T47 + T46;
  assign T46 = nnTop_io_yout_2;
  assign T47 = T48;
  assign T48 = T49;
  assign T49 = T51 + T50;
  assign T50 = nnTop_io_yout_1;
  assign T51 = nnTop_io_yout_0;
  assign io_xout = nnxout;
  assign T52 = T53;
  assign T53 = T55 + T54;
  assign T54 = nnTop_io_xout_2;
  assign T55 = T56;
  assign T56 = T57;
  assign T57 = T59 + T58;
  assign T58 = nnTop_io_xout_1;
  assign T59 = nnTop_io_xout_0;
  NN1Top nnTop(.clk(clk),
       .io_x_2( io_x ),
       .io_x_1( xShift_1 ),
       .io_x_0( xShift_0 ),
       .io_y_11( io_y ),
       .io_y_10( yShift_10 ),
       .io_y_9( yShift_9 ),
       .io_y_8( yShift_8 ),
       .io_y_7( yShift_7 ),
       .io_y_6( yShift_6 ),
       .io_y_5( yShift_5 ),
       .io_y_4( yShift_4 ),
       .io_y_3( yShift_3 ),
       .io_y_2( yShift_2 ),
       .io_y_1( yShift_1 ),
       .io_y_0( yShift_0 ),
       .io_z_2( io_z ),
       .io_z_1( zShift_1 ),
       .io_z_0( zShift_0 ),
       .io_b_11( io_b ),
       .io_b_10( bShift_10 ),
       .io_b_9( bShift_9 ),
       .io_b_8( bShift_8 ),
       .io_b_7( bShift_7 ),
       .io_b_6( bShift_6 ),
       .io_b_5( bShift_5 ),
       .io_b_4( bShift_4 ),
       .io_b_3( bShift_3 ),
       .io_b_2( bShift_2 ),
       .io_b_1( bShift_1 ),
       .io_b_0( bShift_0 ),
       .io_a_11_2( io_a ),
       .io_a_11_1( io_a ),
       .io_a_11_0( io_a ),
       .io_a_10_2( aShift_10_2 ),
       .io_a_10_1( aShift_10_1 ),
       .io_a_10_0( aShift_10_0 ),
       .io_a_9_2( aShift_9_2 ),
       .io_a_9_1( aShift_9_1 ),
       .io_a_9_0( aShift_9_0 ),
       .io_a_8_2( aShift_8_2 ),
       .io_a_8_1( aShift_8_1 ),
       .io_a_8_0( aShift_8_0 ),
       .io_a_7_2( aShift_7_2 ),
       .io_a_7_1( aShift_7_1 ),
       .io_a_7_0( aShift_7_0 ),
       .io_a_6_2( aShift_6_2 ),
       .io_a_6_1( aShift_6_1 ),
       .io_a_6_0( aShift_6_0 ),
       .io_a_5_2( aShift_5_2 ),
       .io_a_5_1( aShift_5_1 ),
       .io_a_5_0( aShift_5_0 ),
       .io_a_4_2( aShift_4_2 ),
       .io_a_4_1( aShift_4_1 ),
       .io_a_4_0( aShift_4_0 ),
       .io_a_3_2( aShift_3_2 ),
       .io_a_3_1( aShift_3_1 ),
       .io_a_3_0( aShift_3_0 ),
       .io_a_2_2( aShift_2_2 ),
       .io_a_2_1( aShift_2_1 ),
       .io_a_2_0( aShift_2_0 ),
       .io_a_1_2( aShift_1_2 ),
       .io_a_1_1( aShift_1_1 ),
       .io_a_1_0( aShift_1_0 ),
       .io_a_0_2( aShift_0_2 ),
       .io_a_0_1( aShift_0_1 ),
       .io_a_0_0( aShift_0_0 ),
       .io_c_2_2( io_c ),
       .io_c_2_1( io_c ),
       .io_c_2_0( io_c ),
       .io_c_1_2( cShift_1_2 ),
       .io_c_1_1( cShift_1_1 ),
       .io_c_1_0( cShift_1_0 ),
       .io_c_0_2( cShift_0_2 ),
       .io_c_0_1( cShift_0_1 ),
       .io_c_0_0( cShift_0_0 ),
       .io_lbda( io_lbda ),
       .io_xout_2( nnTop_io_xout_2 ),
       .io_xout_1( nnTop_io_xout_1 ),
       .io_xout_0( nnTop_io_xout_0 ),
       .io_yout_11( nnTop_io_yout_11 ),
       .io_yout_10( nnTop_io_yout_10 ),
       .io_yout_9( nnTop_io_yout_9 ),
       .io_yout_8( nnTop_io_yout_8 ),
       .io_yout_7( nnTop_io_yout_7 ),
       .io_yout_6( nnTop_io_yout_6 ),
       .io_yout_5( nnTop_io_yout_5 ),
       .io_yout_4( nnTop_io_yout_4 ),
       .io_yout_3( nnTop_io_yout_3 ),
       .io_yout_2( nnTop_io_yout_2 ),
       .io_yout_1( nnTop_io_yout_1 ),
       .io_yout_0( nnTop_io_yout_0 ),
       .io_zout_2( nnTop_io_zout_2 ),
       .io_zout_1( nnTop_io_zout_1 ),
       .io_zout_0( nnTop_io_zout_0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      cShift_0_0 <= 18'h0;
    end else begin
      cShift_0_0 <= cShift_1_0;
    end
    if(reset) begin
      cShift_1_0 <= 18'h0;
    end else begin
      cShift_1_0 <= cShift_2_0;
    end
    if(reset) begin
      cShift_2_0 <= 18'h0;
    end else begin
      cShift_2_0 <= io_c;
    end
    if(reset) begin
      cShift_0_1 <= 18'h0;
    end else begin
      cShift_0_1 <= cShift_1_1;
    end
    if(reset) begin
      cShift_1_1 <= 18'h0;
    end else begin
      cShift_1_1 <= cShift_2_1;
    end
    if(reset) begin
      cShift_2_1 <= 18'h0;
    end else begin
      cShift_2_1 <= io_c;
    end
    if(reset) begin
      cShift_0_2 <= 18'h0;
    end else begin
      cShift_0_2 <= cShift_1_2;
    end
    if(reset) begin
      cShift_1_2 <= 18'h0;
    end else begin
      cShift_1_2 <= cShift_2_2;
    end
    if(reset) begin
      cShift_2_2 <= 18'h0;
    end else begin
      cShift_2_2 <= io_c;
    end
    if(reset) begin
      aShift_0_0 <= 18'h0;
    end else begin
      aShift_0_0 <= aShift_1_0;
    end
    if(reset) begin
      aShift_1_0 <= 18'h0;
    end else begin
      aShift_1_0 <= aShift_2_0;
    end
    if(reset) begin
      aShift_2_0 <= 18'h0;
    end else begin
      aShift_2_0 <= aShift_3_0;
    end
    if(reset) begin
      aShift_3_0 <= 18'h0;
    end else begin
      aShift_3_0 <= aShift_4_0;
    end
    if(reset) begin
      aShift_4_0 <= 18'h0;
    end else begin
      aShift_4_0 <= aShift_5_0;
    end
    if(reset) begin
      aShift_5_0 <= 18'h0;
    end else begin
      aShift_5_0 <= aShift_6_0;
    end
    if(reset) begin
      aShift_6_0 <= 18'h0;
    end else begin
      aShift_6_0 <= aShift_7_0;
    end
    if(reset) begin
      aShift_7_0 <= 18'h0;
    end else begin
      aShift_7_0 <= aShift_8_0;
    end
    if(reset) begin
      aShift_8_0 <= 18'h0;
    end else begin
      aShift_8_0 <= aShift_9_0;
    end
    if(reset) begin
      aShift_9_0 <= 18'h0;
    end else begin
      aShift_9_0 <= aShift_10_0;
    end
    if(reset) begin
      aShift_10_0 <= 18'h0;
    end else begin
      aShift_10_0 <= aShift_11_0;
    end
    if(reset) begin
      aShift_11_0 <= 18'h0;
    end else begin
      aShift_11_0 <= io_a;
    end
    if(reset) begin
      aShift_0_1 <= 18'h0;
    end else begin
      aShift_0_1 <= aShift_1_1;
    end
    if(reset) begin
      aShift_1_1 <= 18'h0;
    end else begin
      aShift_1_1 <= aShift_2_1;
    end
    if(reset) begin
      aShift_2_1 <= 18'h0;
    end else begin
      aShift_2_1 <= aShift_3_1;
    end
    if(reset) begin
      aShift_3_1 <= 18'h0;
    end else begin
      aShift_3_1 <= aShift_4_1;
    end
    if(reset) begin
      aShift_4_1 <= 18'h0;
    end else begin
      aShift_4_1 <= aShift_5_1;
    end
    if(reset) begin
      aShift_5_1 <= 18'h0;
    end else begin
      aShift_5_1 <= aShift_6_1;
    end
    if(reset) begin
      aShift_6_1 <= 18'h0;
    end else begin
      aShift_6_1 <= aShift_7_1;
    end
    if(reset) begin
      aShift_7_1 <= 18'h0;
    end else begin
      aShift_7_1 <= aShift_8_1;
    end
    if(reset) begin
      aShift_8_1 <= 18'h0;
    end else begin
      aShift_8_1 <= aShift_9_1;
    end
    if(reset) begin
      aShift_9_1 <= 18'h0;
    end else begin
      aShift_9_1 <= aShift_10_1;
    end
    if(reset) begin
      aShift_10_1 <= 18'h0;
    end else begin
      aShift_10_1 <= aShift_11_1;
    end
    if(reset) begin
      aShift_11_1 <= 18'h0;
    end else begin
      aShift_11_1 <= io_a;
    end
    if(reset) begin
      aShift_0_2 <= 18'h0;
    end else begin
      aShift_0_2 <= aShift_1_2;
    end
    if(reset) begin
      aShift_1_2 <= 18'h0;
    end else begin
      aShift_1_2 <= aShift_2_2;
    end
    if(reset) begin
      aShift_2_2 <= 18'h0;
    end else begin
      aShift_2_2 <= aShift_3_2;
    end
    if(reset) begin
      aShift_3_2 <= 18'h0;
    end else begin
      aShift_3_2 <= aShift_4_2;
    end
    if(reset) begin
      aShift_4_2 <= 18'h0;
    end else begin
      aShift_4_2 <= aShift_5_2;
    end
    if(reset) begin
      aShift_5_2 <= 18'h0;
    end else begin
      aShift_5_2 <= aShift_6_2;
    end
    if(reset) begin
      aShift_6_2 <= 18'h0;
    end else begin
      aShift_6_2 <= aShift_7_2;
    end
    if(reset) begin
      aShift_7_2 <= 18'h0;
    end else begin
      aShift_7_2 <= aShift_8_2;
    end
    if(reset) begin
      aShift_8_2 <= 18'h0;
    end else begin
      aShift_8_2 <= aShift_9_2;
    end
    if(reset) begin
      aShift_9_2 <= 18'h0;
    end else begin
      aShift_9_2 <= aShift_10_2;
    end
    if(reset) begin
      aShift_10_2 <= 18'h0;
    end else begin
      aShift_10_2 <= aShift_11_2;
    end
    if(reset) begin
      aShift_11_2 <= 18'h0;
    end else begin
      aShift_11_2 <= io_a;
    end
    if(reset) begin
      bShift_0 <= 18'h0;
    end else begin
      bShift_0 <= bShift_1;
    end
    if(reset) begin
      bShift_1 <= 18'h0;
    end else begin
      bShift_1 <= bShift_2;
    end
    if(reset) begin
      bShift_2 <= 18'h0;
    end else begin
      bShift_2 <= bShift_3;
    end
    if(reset) begin
      bShift_3 <= 18'h0;
    end else begin
      bShift_3 <= bShift_4;
    end
    if(reset) begin
      bShift_4 <= 18'h0;
    end else begin
      bShift_4 <= bShift_5;
    end
    if(reset) begin
      bShift_5 <= 18'h0;
    end else begin
      bShift_5 <= bShift_6;
    end
    if(reset) begin
      bShift_6 <= 18'h0;
    end else begin
      bShift_6 <= bShift_7;
    end
    if(reset) begin
      bShift_7 <= 18'h0;
    end else begin
      bShift_7 <= bShift_8;
    end
    if(reset) begin
      bShift_8 <= 18'h0;
    end else begin
      bShift_8 <= bShift_9;
    end
    if(reset) begin
      bShift_9 <= 18'h0;
    end else begin
      bShift_9 <= bShift_10;
    end
    if(reset) begin
      bShift_10 <= 18'h0;
    end else begin
      bShift_10 <= bShift_11;
    end
    if(reset) begin
      bShift_11 <= 18'h0;
    end else begin
      bShift_11 <= io_b;
    end
    if(reset) begin
      zShift_0 <= 18'h0;
    end else begin
      zShift_0 <= zShift_1;
    end
    if(reset) begin
      zShift_1 <= 18'h0;
    end else begin
      zShift_1 <= zShift_2;
    end
    if(reset) begin
      zShift_2 <= 18'h0;
    end else begin
      zShift_2 <= io_z;
    end
    if(reset) begin
      yShift_0 <= 18'h0;
    end else begin
      yShift_0 <= yShift_1;
    end
    if(reset) begin
      yShift_1 <= 18'h0;
    end else begin
      yShift_1 <= yShift_2;
    end
    if(reset) begin
      yShift_2 <= 18'h0;
    end else begin
      yShift_2 <= yShift_3;
    end
    if(reset) begin
      yShift_3 <= 18'h0;
    end else begin
      yShift_3 <= yShift_4;
    end
    if(reset) begin
      yShift_4 <= 18'h0;
    end else begin
      yShift_4 <= yShift_5;
    end
    if(reset) begin
      yShift_5 <= 18'h0;
    end else begin
      yShift_5 <= yShift_6;
    end
    if(reset) begin
      yShift_6 <= 18'h0;
    end else begin
      yShift_6 <= yShift_7;
    end
    if(reset) begin
      yShift_7 <= 18'h0;
    end else begin
      yShift_7 <= yShift_8;
    end
    if(reset) begin
      yShift_8 <= 18'h0;
    end else begin
      yShift_8 <= yShift_9;
    end
    if(reset) begin
      yShift_9 <= 18'h0;
    end else begin
      yShift_9 <= yShift_10;
    end
    if(reset) begin
      yShift_10 <= 18'h0;
    end else begin
      yShift_10 <= yShift_11;
    end
    if(reset) begin
      yShift_11 <= 18'h0;
    end else begin
      yShift_11 <= io_y;
    end
    if(reset) begin
      xShift_0 <= 18'h0;
    end else begin
      xShift_0 <= xShift_1;
    end
    if(reset) begin
      xShift_1 <= 18'h0;
    end else begin
      xShift_1 <= xShift_2;
    end
    if(reset) begin
      xShift_2 <= 18'h0;
    end else begin
      xShift_2 <= io_x;
    end
    nnzout <= T0;
    nnyout <= T8;
    nnxout <= T52;
  end
endmodule

