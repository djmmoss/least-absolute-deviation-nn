module XNetModule(
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_y_11,
    input [17:0] io_y_10,
    input [17:0] io_y_9,
    input [17:0] io_y_8,
    input [17:0] io_y_7,
    input [17:0] io_y_6,
    input [17:0] io_y_5,
    input [17:0] io_y_4,
    input [17:0] io_y_3,
    input [17:0] io_y_2,
    input [17:0] io_y_1,
    input [17:0] io_y_0,
    input [17:0] io_z_2,
    input [17:0] io_z_1,
    input [17:0] io_z_0,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_c_2_2,
    input [17:0] io_c_2_1,
    input [17:0] io_c_2_0,
    input [17:0] io_c_1_2,
    input [17:0] io_c_1_1,
    input [17:0] io_c_1_0,
    input [17:0] io_c_0_2,
    input [17:0] io_c_0_1,
    input [17:0] io_c_0_0,
    output[17:0] io_o_2,
    output[17:0] io_o_1,
    output[17:0] io_o_0
);

  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] x_stage_0;
  wire[17:0] T2;
  wire[17:0] T3;
  wire[17:0] cz_0;
  wire[17:0] T4;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T417;
  wire[21:0] T7;
  wire[35:0] T8;
  wire[17:0] T9;
  wire[17:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  wire[17:0] T418;
  wire[21:0] T16;
  wire[35:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  wire[17:0] T20;
  wire[17:0] T21;
  wire[17:0] T419;
  wire[21:0] T22;
  wire[35:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;
  wire[17:0] T26;
  wire[17:0] xay_0;
  wire[17:0] T27;
  wire[17:0] T28;
  wire[17:0] ay_0;
  wire[17:0] T29;
  wire[17:0] T30;
  wire[17:0] T31;
  wire[17:0] T32;
  wire[17:0] T33;
  wire[17:0] T34;
  wire[17:0] T35;
  wire[17:0] T36;
  wire[17:0] T37;
  wire[17:0] T420;
  wire[21:0] T38;
  wire[35:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  wire[17:0] T42;
  wire[17:0] T43;
  wire[17:0] T421;
  wire[21:0] T44;
  wire[35:0] T45;
  wire[17:0] T46;
  wire[17:0] T47;
  wire[17:0] T48;
  wire[17:0] T49;
  wire[17:0] T50;
  wire[17:0] T51;
  wire[17:0] T52;
  wire[17:0] T422;
  wire[21:0] T53;
  wire[35:0] T54;
  wire[17:0] T55;
  wire[17:0] T56;
  wire[17:0] T57;
  wire[17:0] T58;
  wire[17:0] T423;
  wire[21:0] T59;
  wire[35:0] T60;
  wire[17:0] T61;
  wire[17:0] T62;
  wire[17:0] T63;
  wire[17:0] T64;
  wire[17:0] T65;
  wire[17:0] T66;
  wire[17:0] T67;
  wire[17:0] T68;
  wire[17:0] T69;
  wire[17:0] T70;
  wire[17:0] T71;
  wire[17:0] T72;
  wire[17:0] T73;
  wire[17:0] T424;
  wire[21:0] T74;
  wire[35:0] T75;
  wire[17:0] T76;
  wire[17:0] T77;
  wire[17:0] T78;
  wire[17:0] T79;
  wire[17:0] T425;
  wire[21:0] T80;
  wire[35:0] T81;
  wire[17:0] T82;
  wire[17:0] T83;
  wire[17:0] T84;
  wire[17:0] T85;
  wire[17:0] T86;
  wire[17:0] T87;
  wire[17:0] T88;
  wire[17:0] T426;
  wire[21:0] T89;
  wire[35:0] T90;
  wire[17:0] T91;
  wire[17:0] T92;
  wire[17:0] T93;
  wire[17:0] T94;
  wire[17:0] T427;
  wire[21:0] T95;
  wire[35:0] T96;
  wire[17:0] T97;
  wire[17:0] T98;
  wire[17:0] T99;
  wire[17:0] T100;
  wire[17:0] T101;
  wire[17:0] T102;
  wire[17:0] T103;
  wire[17:0] T104;
  wire[17:0] T105;
  wire[17:0] T106;
  wire[17:0] T428;
  wire[21:0] T107;
  wire[35:0] T108;
  wire[17:0] T109;
  wire[17:0] T110;
  wire[17:0] T111;
  wire[17:0] T112;
  wire[17:0] T429;
  wire[21:0] T113;
  wire[35:0] T114;
  wire[17:0] T115;
  wire[17:0] T116;
  wire[17:0] T117;
  wire[17:0] T118;
  wire[17:0] T119;
  wire[17:0] T120;
  wire[17:0] T121;
  wire[17:0] T430;
  wire[21:0] T122;
  wire[35:0] T123;
  wire[17:0] T124;
  wire[17:0] T125;
  wire[17:0] T126;
  wire[17:0] T127;
  wire[17:0] T431;
  wire[21:0] T128;
  wire[35:0] T129;
  wire[17:0] T130;
  wire[17:0] T131;
  wire[17:0] T132;
  wire T133;
  wire[17:0] T134;
  wire[17:0] T135;
  wire T136;
  wire[17:0] T137;
  wire[17:0] T138;
  wire[17:0] T139;
  wire[17:0] T140;
  wire[17:0] x_stage_1;
  wire[17:0] T141;
  wire[17:0] T142;
  wire[17:0] cz_1;
  wire[17:0] T143;
  wire[17:0] T144;
  wire[17:0] T145;
  wire[17:0] T432;
  wire[21:0] T146;
  wire[35:0] T147;
  wire[17:0] T148;
  wire[17:0] T149;
  wire[17:0] T150;
  wire[17:0] T151;
  wire[17:0] T152;
  wire[17:0] T153;
  wire[17:0] T154;
  wire[17:0] T433;
  wire[21:0] T155;
  wire[35:0] T156;
  wire[17:0] T157;
  wire[17:0] T158;
  wire[17:0] T159;
  wire[17:0] T160;
  wire[17:0] T434;
  wire[21:0] T161;
  wire[35:0] T162;
  wire[17:0] T163;
  wire[17:0] T164;
  wire[17:0] T165;
  wire[17:0] xay_1;
  wire[17:0] T166;
  wire[17:0] T167;
  wire[17:0] ay_1;
  wire[17:0] T168;
  wire[17:0] T169;
  wire[17:0] T170;
  wire[17:0] T171;
  wire[17:0] T172;
  wire[17:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[17:0] T176;
  wire[17:0] T435;
  wire[21:0] T177;
  wire[35:0] T178;
  wire[17:0] T179;
  wire[17:0] T180;
  wire[17:0] T181;
  wire[17:0] T182;
  wire[17:0] T436;
  wire[21:0] T183;
  wire[35:0] T184;
  wire[17:0] T185;
  wire[17:0] T186;
  wire[17:0] T187;
  wire[17:0] T188;
  wire[17:0] T189;
  wire[17:0] T190;
  wire[17:0] T191;
  wire[17:0] T437;
  wire[21:0] T192;
  wire[35:0] T193;
  wire[17:0] T194;
  wire[17:0] T195;
  wire[17:0] T196;
  wire[17:0] T197;
  wire[17:0] T438;
  wire[21:0] T198;
  wire[35:0] T199;
  wire[17:0] T200;
  wire[17:0] T201;
  wire[17:0] T202;
  wire[17:0] T203;
  wire[17:0] T204;
  wire[17:0] T205;
  wire[17:0] T206;
  wire[17:0] T207;
  wire[17:0] T208;
  wire[17:0] T209;
  wire[17:0] T210;
  wire[17:0] T211;
  wire[17:0] T212;
  wire[17:0] T439;
  wire[21:0] T213;
  wire[35:0] T214;
  wire[17:0] T215;
  wire[17:0] T216;
  wire[17:0] T217;
  wire[17:0] T218;
  wire[17:0] T440;
  wire[21:0] T219;
  wire[35:0] T220;
  wire[17:0] T221;
  wire[17:0] T222;
  wire[17:0] T223;
  wire[17:0] T224;
  wire[17:0] T225;
  wire[17:0] T226;
  wire[17:0] T227;
  wire[17:0] T441;
  wire[21:0] T228;
  wire[35:0] T229;
  wire[17:0] T230;
  wire[17:0] T231;
  wire[17:0] T232;
  wire[17:0] T233;
  wire[17:0] T442;
  wire[21:0] T234;
  wire[35:0] T235;
  wire[17:0] T236;
  wire[17:0] T237;
  wire[17:0] T238;
  wire[17:0] T239;
  wire[17:0] T240;
  wire[17:0] T241;
  wire[17:0] T242;
  wire[17:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[17:0] T443;
  wire[21:0] T246;
  wire[35:0] T247;
  wire[17:0] T248;
  wire[17:0] T249;
  wire[17:0] T250;
  wire[17:0] T251;
  wire[17:0] T444;
  wire[21:0] T252;
  wire[35:0] T253;
  wire[17:0] T254;
  wire[17:0] T255;
  wire[17:0] T256;
  wire[17:0] T257;
  wire[17:0] T258;
  wire[17:0] T259;
  wire[17:0] T260;
  wire[17:0] T445;
  wire[21:0] T261;
  wire[35:0] T262;
  wire[17:0] T263;
  wire[17:0] T264;
  wire[17:0] T265;
  wire[17:0] T266;
  wire[17:0] T446;
  wire[21:0] T267;
  wire[35:0] T268;
  wire[17:0] T269;
  wire[17:0] T270;
  wire[17:0] T271;
  wire T272;
  wire[17:0] T273;
  wire[17:0] T274;
  wire T275;
  wire[17:0] T276;
  wire[17:0] T277;
  wire[17:0] T278;
  wire[17:0] T279;
  wire[17:0] x_stage_2;
  wire[17:0] T280;
  wire[17:0] T281;
  wire[17:0] cz_2;
  wire[17:0] T282;
  wire[17:0] T283;
  wire[17:0] T284;
  wire[17:0] T447;
  wire[21:0] T285;
  wire[35:0] T286;
  wire[17:0] T287;
  wire[17:0] T288;
  wire[17:0] T289;
  wire[17:0] T290;
  wire[17:0] T291;
  wire[17:0] T292;
  wire[17:0] T293;
  wire[17:0] T448;
  wire[21:0] T294;
  wire[35:0] T295;
  wire[17:0] T296;
  wire[17:0] T297;
  wire[17:0] T298;
  wire[17:0] T299;
  wire[17:0] T449;
  wire[21:0] T300;
  wire[35:0] T301;
  wire[17:0] T302;
  wire[17:0] T303;
  wire[17:0] T304;
  wire[17:0] xay_2;
  wire[17:0] T305;
  wire[17:0] T306;
  wire[17:0] ay_2;
  wire[17:0] T307;
  wire[17:0] T308;
  wire[17:0] T309;
  wire[17:0] T310;
  wire[17:0] T311;
  wire[17:0] T312;
  wire[17:0] T313;
  wire[17:0] T314;
  wire[17:0] T315;
  wire[17:0] T450;
  wire[21:0] T316;
  wire[35:0] T317;
  wire[17:0] T318;
  wire[17:0] T319;
  wire[17:0] T320;
  wire[17:0] T321;
  wire[17:0] T451;
  wire[21:0] T322;
  wire[35:0] T323;
  wire[17:0] T324;
  wire[17:0] T325;
  wire[17:0] T326;
  wire[17:0] T327;
  wire[17:0] T328;
  wire[17:0] T329;
  wire[17:0] T330;
  wire[17:0] T452;
  wire[21:0] T331;
  wire[35:0] T332;
  wire[17:0] T333;
  wire[17:0] T334;
  wire[17:0] T335;
  wire[17:0] T336;
  wire[17:0] T453;
  wire[21:0] T337;
  wire[35:0] T338;
  wire[17:0] T339;
  wire[17:0] T340;
  wire[17:0] T341;
  wire[17:0] T342;
  wire[17:0] T343;
  wire[17:0] T344;
  wire[17:0] T345;
  wire[17:0] T346;
  wire[17:0] T347;
  wire[17:0] T348;
  wire[17:0] T349;
  wire[17:0] T350;
  wire[17:0] T351;
  wire[17:0] T454;
  wire[21:0] T352;
  wire[35:0] T353;
  wire[17:0] T354;
  wire[17:0] T355;
  wire[17:0] T356;
  wire[17:0] T357;
  wire[17:0] T455;
  wire[21:0] T358;
  wire[35:0] T359;
  wire[17:0] T360;
  wire[17:0] T361;
  wire[17:0] T362;
  wire[17:0] T363;
  wire[17:0] T364;
  wire[17:0] T365;
  wire[17:0] T366;
  wire[17:0] T456;
  wire[21:0] T367;
  wire[35:0] T368;
  wire[17:0] T369;
  wire[17:0] T370;
  wire[17:0] T371;
  wire[17:0] T372;
  wire[17:0] T457;
  wire[21:0] T373;
  wire[35:0] T374;
  wire[17:0] T375;
  wire[17:0] T376;
  wire[17:0] T377;
  wire[17:0] T378;
  wire[17:0] T379;
  wire[17:0] T380;
  wire[17:0] T381;
  wire[17:0] T382;
  wire[17:0] T383;
  wire[17:0] T384;
  wire[17:0] T458;
  wire[21:0] T385;
  wire[35:0] T386;
  wire[17:0] T387;
  wire[17:0] T388;
  wire[17:0] T389;
  wire[17:0] T390;
  wire[17:0] T459;
  wire[21:0] T391;
  wire[35:0] T392;
  wire[17:0] T393;
  wire[17:0] T394;
  wire[17:0] T395;
  wire[17:0] T396;
  wire[17:0] T397;
  wire[17:0] T398;
  wire[17:0] T399;
  wire[17:0] T460;
  wire[21:0] T400;
  wire[35:0] T401;
  wire[17:0] T402;
  wire[17:0] T403;
  wire[17:0] T404;
  wire[17:0] T405;
  wire[17:0] T461;
  wire[21:0] T406;
  wire[35:0] T407;
  wire[17:0] T408;
  wire[17:0] T409;
  wire[17:0] T410;
  wire T411;
  wire[17:0] T412;
  wire[17:0] T413;
  wire T414;
  wire[17:0] T415;
  wire[17:0] T416;


  assign io_o_0 = T0;
  assign T0 = T136 ? 18'h8000 : T1;
  assign T1 = T133 ? 18'h38000 : x_stage_0;
  assign x_stage_0 = T2;
  assign T2 = T26 + T3;
  assign T3 = cz_0;
  assign cz_0 = T4;
  assign T4 = T11 + T5;
  assign T5 = T6;
  assign T6 = T417;
  assign T417 = T7[5'h11:1'h0];
  assign T7 = $signed(T8) >>> 4'he;
  assign T8 = $signed(T10) * $signed(T9);
  assign T9 = io_z_2;
  assign T10 = io_c_2_0;
  assign T11 = T12;
  assign T12 = T13;
  assign T13 = T20 + T14;
  assign T14 = T15;
  assign T15 = T418;
  assign T418 = T16[5'h11:1'h0];
  assign T16 = $signed(T17) >>> 4'he;
  assign T17 = $signed(T19) * $signed(T18);
  assign T18 = io_z_1;
  assign T19 = io_c_1_0;
  assign T20 = T21;
  assign T21 = T419;
  assign T419 = T22[5'h11:1'h0];
  assign T22 = $signed(T23) >>> 4'he;
  assign T23 = $signed(T25) * $signed(T24);
  assign T24 = io_z_0;
  assign T25 = io_c_0_0;
  assign T26 = xay_0;
  assign xay_0 = T27;
  assign T27 = T132 - T28;
  assign T28 = ay_0;
  assign ay_0 = T29;
  assign T29 = T63 + T30;
  assign T30 = T31;
  assign T31 = T32;
  assign T32 = T48 + T33;
  assign T33 = T34;
  assign T34 = T35;
  assign T35 = T42 + T36;
  assign T36 = T37;
  assign T37 = T420;
  assign T420 = T38[5'h11:1'h0];
  assign T38 = $signed(T39) >>> 4'he;
  assign T39 = $signed(T41) * $signed(T40);
  assign T40 = io_y_11;
  assign T41 = io_a_11_0;
  assign T42 = T43;
  assign T43 = T421;
  assign T421 = T44[5'h11:1'h0];
  assign T44 = $signed(T45) >>> 4'he;
  assign T45 = $signed(T47) * $signed(T46);
  assign T46 = io_y_10;
  assign T47 = io_a_10_0;
  assign T48 = T49;
  assign T49 = T50;
  assign T50 = T57 + T51;
  assign T51 = T52;
  assign T52 = T422;
  assign T422 = T53[5'h11:1'h0];
  assign T53 = $signed(T54) >>> 4'he;
  assign T54 = $signed(T56) * $signed(T55);
  assign T55 = io_y_9;
  assign T56 = io_a_9_0;
  assign T57 = T58;
  assign T58 = T423;
  assign T423 = T59[5'h11:1'h0];
  assign T59 = $signed(T60) >>> 4'he;
  assign T60 = $signed(T62) * $signed(T61);
  assign T61 = io_y_8;
  assign T62 = io_a_8_0;
  assign T63 = T64;
  assign T64 = T65;
  assign T65 = T99 + T66;
  assign T66 = T67;
  assign T67 = T68;
  assign T68 = T84 + T69;
  assign T69 = T70;
  assign T70 = T71;
  assign T71 = T78 + T72;
  assign T72 = T73;
  assign T73 = T424;
  assign T424 = T74[5'h11:1'h0];
  assign T74 = $signed(T75) >>> 4'he;
  assign T75 = $signed(T77) * $signed(T76);
  assign T76 = io_y_7;
  assign T77 = io_a_7_0;
  assign T78 = T79;
  assign T79 = T425;
  assign T425 = T80[5'h11:1'h0];
  assign T80 = $signed(T81) >>> 4'he;
  assign T81 = $signed(T83) * $signed(T82);
  assign T82 = io_y_6;
  assign T83 = io_a_6_0;
  assign T84 = T85;
  assign T85 = T86;
  assign T86 = T93 + T87;
  assign T87 = T88;
  assign T88 = T426;
  assign T426 = T89[5'h11:1'h0];
  assign T89 = $signed(T90) >>> 4'he;
  assign T90 = $signed(T92) * $signed(T91);
  assign T91 = io_y_5;
  assign T92 = io_a_5_0;
  assign T93 = T94;
  assign T94 = T427;
  assign T427 = T95[5'h11:1'h0];
  assign T95 = $signed(T96) >>> 4'he;
  assign T96 = $signed(T98) * $signed(T97);
  assign T97 = io_y_4;
  assign T98 = io_a_4_0;
  assign T99 = T100;
  assign T100 = T101;
  assign T101 = T117 + T102;
  assign T102 = T103;
  assign T103 = T104;
  assign T104 = T111 + T105;
  assign T105 = T106;
  assign T106 = T428;
  assign T428 = T107[5'h11:1'h0];
  assign T107 = $signed(T108) >>> 4'he;
  assign T108 = $signed(T110) * $signed(T109);
  assign T109 = io_y_3;
  assign T110 = io_a_3_0;
  assign T111 = T112;
  assign T112 = T429;
  assign T429 = T113[5'h11:1'h0];
  assign T113 = $signed(T114) >>> 4'he;
  assign T114 = $signed(T116) * $signed(T115);
  assign T115 = io_y_2;
  assign T116 = io_a_2_0;
  assign T117 = T118;
  assign T118 = T119;
  assign T119 = T126 + T120;
  assign T120 = T121;
  assign T121 = T430;
  assign T430 = T122[5'h11:1'h0];
  assign T122 = $signed(T123) >>> 4'he;
  assign T123 = $signed(T125) * $signed(T124);
  assign T124 = io_y_1;
  assign T125 = io_a_1_0;
  assign T126 = T127;
  assign T127 = T431;
  assign T431 = T128[5'h11:1'h0];
  assign T128 = $signed(T129) >>> 4'he;
  assign T129 = $signed(T131) * $signed(T130);
  assign T130 = io_y_0;
  assign T131 = io_a_0_0;
  assign T132 = io_x_0;
  assign T133 = $signed(T135) < $signed(T134);
  assign T134 = 18'h38000;
  assign T135 = x_stage_0;
  assign T136 = $signed(T138) < $signed(T137);
  assign T137 = x_stage_0;
  assign T138 = 18'h8000;
  assign io_o_1 = T139;
  assign T139 = T275 ? 18'h8000 : T140;
  assign T140 = T272 ? 18'h38000 : x_stage_1;
  assign x_stage_1 = T141;
  assign T141 = T165 + T142;
  assign T142 = cz_1;
  assign cz_1 = T143;
  assign T143 = T150 + T144;
  assign T144 = T145;
  assign T145 = T432;
  assign T432 = T146[5'h11:1'h0];
  assign T146 = $signed(T147) >>> 4'he;
  assign T147 = $signed(T149) * $signed(T148);
  assign T148 = io_z_2;
  assign T149 = io_c_2_1;
  assign T150 = T151;
  assign T151 = T152;
  assign T152 = T159 + T153;
  assign T153 = T154;
  assign T154 = T433;
  assign T433 = T155[5'h11:1'h0];
  assign T155 = $signed(T156) >>> 4'he;
  assign T156 = $signed(T158) * $signed(T157);
  assign T157 = io_z_1;
  assign T158 = io_c_1_1;
  assign T159 = T160;
  assign T160 = T434;
  assign T434 = T161[5'h11:1'h0];
  assign T161 = $signed(T162) >>> 4'he;
  assign T162 = $signed(T164) * $signed(T163);
  assign T163 = io_z_0;
  assign T164 = io_c_0_1;
  assign T165 = xay_1;
  assign xay_1 = T166;
  assign T166 = T271 - T167;
  assign T167 = ay_1;
  assign ay_1 = T168;
  assign T168 = T202 + T169;
  assign T169 = T170;
  assign T170 = T171;
  assign T171 = T187 + T172;
  assign T172 = T173;
  assign T173 = T174;
  assign T174 = T181 + T175;
  assign T175 = T176;
  assign T176 = T435;
  assign T435 = T177[5'h11:1'h0];
  assign T177 = $signed(T178) >>> 4'he;
  assign T178 = $signed(T180) * $signed(T179);
  assign T179 = io_y_11;
  assign T180 = io_a_11_1;
  assign T181 = T182;
  assign T182 = T436;
  assign T436 = T183[5'h11:1'h0];
  assign T183 = $signed(T184) >>> 4'he;
  assign T184 = $signed(T186) * $signed(T185);
  assign T185 = io_y_10;
  assign T186 = io_a_10_1;
  assign T187 = T188;
  assign T188 = T189;
  assign T189 = T196 + T190;
  assign T190 = T191;
  assign T191 = T437;
  assign T437 = T192[5'h11:1'h0];
  assign T192 = $signed(T193) >>> 4'he;
  assign T193 = $signed(T195) * $signed(T194);
  assign T194 = io_y_9;
  assign T195 = io_a_9_1;
  assign T196 = T197;
  assign T197 = T438;
  assign T438 = T198[5'h11:1'h0];
  assign T198 = $signed(T199) >>> 4'he;
  assign T199 = $signed(T201) * $signed(T200);
  assign T200 = io_y_8;
  assign T201 = io_a_8_1;
  assign T202 = T203;
  assign T203 = T204;
  assign T204 = T238 + T205;
  assign T205 = T206;
  assign T206 = T207;
  assign T207 = T223 + T208;
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T217 + T211;
  assign T211 = T212;
  assign T212 = T439;
  assign T439 = T213[5'h11:1'h0];
  assign T213 = $signed(T214) >>> 4'he;
  assign T214 = $signed(T216) * $signed(T215);
  assign T215 = io_y_7;
  assign T216 = io_a_7_1;
  assign T217 = T218;
  assign T218 = T440;
  assign T440 = T219[5'h11:1'h0];
  assign T219 = $signed(T220) >>> 4'he;
  assign T220 = $signed(T222) * $signed(T221);
  assign T221 = io_y_6;
  assign T222 = io_a_6_1;
  assign T223 = T224;
  assign T224 = T225;
  assign T225 = T232 + T226;
  assign T226 = T227;
  assign T227 = T441;
  assign T441 = T228[5'h11:1'h0];
  assign T228 = $signed(T229) >>> 4'he;
  assign T229 = $signed(T231) * $signed(T230);
  assign T230 = io_y_5;
  assign T231 = io_a_5_1;
  assign T232 = T233;
  assign T233 = T442;
  assign T442 = T234[5'h11:1'h0];
  assign T234 = $signed(T235) >>> 4'he;
  assign T235 = $signed(T237) * $signed(T236);
  assign T236 = io_y_4;
  assign T237 = io_a_4_1;
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T256 + T241;
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = T250 + T244;
  assign T244 = T245;
  assign T245 = T443;
  assign T443 = T246[5'h11:1'h0];
  assign T246 = $signed(T247) >>> 4'he;
  assign T247 = $signed(T249) * $signed(T248);
  assign T248 = io_y_3;
  assign T249 = io_a_3_1;
  assign T250 = T251;
  assign T251 = T444;
  assign T444 = T252[5'h11:1'h0];
  assign T252 = $signed(T253) >>> 4'he;
  assign T253 = $signed(T255) * $signed(T254);
  assign T254 = io_y_2;
  assign T255 = io_a_2_1;
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T265 + T259;
  assign T259 = T260;
  assign T260 = T445;
  assign T445 = T261[5'h11:1'h0];
  assign T261 = $signed(T262) >>> 4'he;
  assign T262 = $signed(T264) * $signed(T263);
  assign T263 = io_y_1;
  assign T264 = io_a_1_1;
  assign T265 = T266;
  assign T266 = T446;
  assign T446 = T267[5'h11:1'h0];
  assign T267 = $signed(T268) >>> 4'he;
  assign T268 = $signed(T270) * $signed(T269);
  assign T269 = io_y_0;
  assign T270 = io_a_0_1;
  assign T271 = io_x_1;
  assign T272 = $signed(T274) < $signed(T273);
  assign T273 = 18'h38000;
  assign T274 = x_stage_1;
  assign T275 = $signed(T277) < $signed(T276);
  assign T276 = x_stage_1;
  assign T277 = 18'h8000;
  assign io_o_2 = T278;
  assign T278 = T414 ? 18'h8000 : T279;
  assign T279 = T411 ? 18'h38000 : x_stage_2;
  assign x_stage_2 = T280;
  assign T280 = T304 + T281;
  assign T281 = cz_2;
  assign cz_2 = T282;
  assign T282 = T289 + T283;
  assign T283 = T284;
  assign T284 = T447;
  assign T447 = T285[5'h11:1'h0];
  assign T285 = $signed(T286) >>> 4'he;
  assign T286 = $signed(T288) * $signed(T287);
  assign T287 = io_z_2;
  assign T288 = io_c_2_2;
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = T298 + T292;
  assign T292 = T293;
  assign T293 = T448;
  assign T448 = T294[5'h11:1'h0];
  assign T294 = $signed(T295) >>> 4'he;
  assign T295 = $signed(T297) * $signed(T296);
  assign T296 = io_z_1;
  assign T297 = io_c_1_2;
  assign T298 = T299;
  assign T299 = T449;
  assign T449 = T300[5'h11:1'h0];
  assign T300 = $signed(T301) >>> 4'he;
  assign T301 = $signed(T303) * $signed(T302);
  assign T302 = io_z_0;
  assign T303 = io_c_0_2;
  assign T304 = xay_2;
  assign xay_2 = T305;
  assign T305 = T410 - T306;
  assign T306 = ay_2;
  assign ay_2 = T307;
  assign T307 = T341 + T308;
  assign T308 = T309;
  assign T309 = T310;
  assign T310 = T326 + T311;
  assign T311 = T312;
  assign T312 = T313;
  assign T313 = T320 + T314;
  assign T314 = T315;
  assign T315 = T450;
  assign T450 = T316[5'h11:1'h0];
  assign T316 = $signed(T317) >>> 4'he;
  assign T317 = $signed(T319) * $signed(T318);
  assign T318 = io_y_11;
  assign T319 = io_a_11_2;
  assign T320 = T321;
  assign T321 = T451;
  assign T451 = T322[5'h11:1'h0];
  assign T322 = $signed(T323) >>> 4'he;
  assign T323 = $signed(T325) * $signed(T324);
  assign T324 = io_y_10;
  assign T325 = io_a_10_2;
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T335 + T329;
  assign T329 = T330;
  assign T330 = T452;
  assign T452 = T331[5'h11:1'h0];
  assign T331 = $signed(T332) >>> 4'he;
  assign T332 = $signed(T334) * $signed(T333);
  assign T333 = io_y_9;
  assign T334 = io_a_9_2;
  assign T335 = T336;
  assign T336 = T453;
  assign T453 = T337[5'h11:1'h0];
  assign T337 = $signed(T338) >>> 4'he;
  assign T338 = $signed(T340) * $signed(T339);
  assign T339 = io_y_8;
  assign T340 = io_a_8_2;
  assign T341 = T342;
  assign T342 = T343;
  assign T343 = T377 + T344;
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T362 + T347;
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = T356 + T350;
  assign T350 = T351;
  assign T351 = T454;
  assign T454 = T352[5'h11:1'h0];
  assign T352 = $signed(T353) >>> 4'he;
  assign T353 = $signed(T355) * $signed(T354);
  assign T354 = io_y_7;
  assign T355 = io_a_7_2;
  assign T356 = T357;
  assign T357 = T455;
  assign T455 = T358[5'h11:1'h0];
  assign T358 = $signed(T359) >>> 4'he;
  assign T359 = $signed(T361) * $signed(T360);
  assign T360 = io_y_6;
  assign T361 = io_a_6_2;
  assign T362 = T363;
  assign T363 = T364;
  assign T364 = T371 + T365;
  assign T365 = T366;
  assign T366 = T456;
  assign T456 = T367[5'h11:1'h0];
  assign T367 = $signed(T368) >>> 4'he;
  assign T368 = $signed(T370) * $signed(T369);
  assign T369 = io_y_5;
  assign T370 = io_a_5_2;
  assign T371 = T372;
  assign T372 = T457;
  assign T457 = T373[5'h11:1'h0];
  assign T373 = $signed(T374) >>> 4'he;
  assign T374 = $signed(T376) * $signed(T375);
  assign T375 = io_y_4;
  assign T376 = io_a_4_2;
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = T395 + T380;
  assign T380 = T381;
  assign T381 = T382;
  assign T382 = T389 + T383;
  assign T383 = T384;
  assign T384 = T458;
  assign T458 = T385[5'h11:1'h0];
  assign T385 = $signed(T386) >>> 4'he;
  assign T386 = $signed(T388) * $signed(T387);
  assign T387 = io_y_3;
  assign T388 = io_a_3_2;
  assign T389 = T390;
  assign T390 = T459;
  assign T459 = T391[5'h11:1'h0];
  assign T391 = $signed(T392) >>> 4'he;
  assign T392 = $signed(T394) * $signed(T393);
  assign T393 = io_y_2;
  assign T394 = io_a_2_2;
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = T404 + T398;
  assign T398 = T399;
  assign T399 = T460;
  assign T460 = T400[5'h11:1'h0];
  assign T400 = $signed(T401) >>> 4'he;
  assign T401 = $signed(T403) * $signed(T402);
  assign T402 = io_y_1;
  assign T403 = io_a_1_2;
  assign T404 = T405;
  assign T405 = T461;
  assign T461 = T406[5'h11:1'h0];
  assign T406 = $signed(T407) >>> 4'he;
  assign T407 = $signed(T409) * $signed(T408);
  assign T408 = io_y_0;
  assign T409 = io_a_0_2;
  assign T410 = io_x_2;
  assign T411 = $signed(T413) < $signed(T412);
  assign T412 = 18'h38000;
  assign T413 = x_stage_2;
  assign T414 = $signed(T416) < $signed(T415);
  assign T415 = x_stage_2;
  assign T416 = 18'h8000;
endmodule

module NN1Top(input clk,
    input [17:0] io_x_2,
    input [17:0] io_x_1,
    input [17:0] io_x_0,
    input [17:0] io_y_11,
    input [17:0] io_y_10,
    input [17:0] io_y_9,
    input [17:0] io_y_8,
    input [17:0] io_y_7,
    input [17:0] io_y_6,
    input [17:0] io_y_5,
    input [17:0] io_y_4,
    input [17:0] io_y_3,
    input [17:0] io_y_2,
    input [17:0] io_y_1,
    input [17:0] io_y_0,
    input [17:0] io_z_2,
    input [17:0] io_z_1,
    input [17:0] io_z_0,
    input [17:0] io_b_11,
    input [17:0] io_b_10,
    input [17:0] io_b_9,
    input [17:0] io_b_8,
    input [17:0] io_b_7,
    input [17:0] io_b_6,
    input [17:0] io_b_5,
    input [17:0] io_b_4,
    input [17:0] io_b_3,
    input [17:0] io_b_2,
    input [17:0] io_b_1,
    input [17:0] io_b_0,
    input [17:0] io_a_11_2,
    input [17:0] io_a_11_1,
    input [17:0] io_a_11_0,
    input [17:0] io_a_10_2,
    input [17:0] io_a_10_1,
    input [17:0] io_a_10_0,
    input [17:0] io_a_9_2,
    input [17:0] io_a_9_1,
    input [17:0] io_a_9_0,
    input [17:0] io_a_8_2,
    input [17:0] io_a_8_1,
    input [17:0] io_a_8_0,
    input [17:0] io_a_7_2,
    input [17:0] io_a_7_1,
    input [17:0] io_a_7_0,
    input [17:0] io_a_6_2,
    input [17:0] io_a_6_1,
    input [17:0] io_a_6_0,
    input [17:0] io_a_5_2,
    input [17:0] io_a_5_1,
    input [17:0] io_a_5_0,
    input [17:0] io_a_4_2,
    input [17:0] io_a_4_1,
    input [17:0] io_a_4_0,
    input [17:0] io_a_3_2,
    input [17:0] io_a_3_1,
    input [17:0] io_a_3_0,
    input [17:0] io_a_2_2,
    input [17:0] io_a_2_1,
    input [17:0] io_a_2_0,
    input [17:0] io_a_1_2,
    input [17:0] io_a_1_1,
    input [17:0] io_a_1_0,
    input [17:0] io_a_0_2,
    input [17:0] io_a_0_1,
    input [17:0] io_a_0_0,
    input [17:0] io_c_2_2,
    input [17:0] io_c_2_1,
    input [17:0] io_c_2_0,
    input [17:0] io_c_1_2,
    input [17:0] io_c_1_1,
    input [17:0] io_c_1_0,
    input [17:0] io_c_0_2,
    input [17:0] io_c_0_1,
    input [17:0] io_c_0_0,
    input [17:0] io_lbda,
    output[17:0] io_xout_2,
    output[17:0] io_xout_1,
    output[17:0] io_xout_0,
    output[17:0] io_yout_11,
    output[17:0] io_yout_10,
    output[17:0] io_yout_9,
    output[17:0] io_yout_8,
    output[17:0] io_yout_7,
    output[17:0] io_yout_6,
    output[17:0] io_yout_5,
    output[17:0] io_yout_4,
    output[17:0] io_yout_3,
    output[17:0] io_yout_2,
    output[17:0] io_yout_1,
    output[17:0] io_yout_0,
    output[17:0] io_zout_2,
    output[17:0] io_zout_1,
    output[17:0] io_zout_0
);

  wire[17:0] zout_0;
  wire[17:0] T0;
  wire[17:0] T1;
  reg [17:0] R2;
  wire[17:0] T3;
  wire[17:0] T1134;
  wire[21:0] T4;
  wire[35:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  wire[17:0] T8;
  wire[17:0] T1135;
  wire[21:0] T9;
  wire[35:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  reg [17:0] R16;
  wire[17:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  wire[17:0] T20;
  wire[17:0] T21;
  reg [17:0] R22;
  reg [17:0] R23;
  wire[17:0] T24;
  wire[17:0] T25;
  wire[17:0] T26;
  wire[17:0] T27;
  wire[17:0] T28;
  wire[17:0] T1136;
  wire[21:0] T29;
  wire[35:0] T30;
  wire[17:0] T31;
  reg [17:0] R32;
  reg [17:0] R33;
  wire[17:0] T34;
  reg [17:0] R35;
  reg [17:0] R36;
  wire[17:0] T37;
  wire[17:0] T38;
  wire[17:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  wire[17:0] T1137;
  wire[21:0] T42;
  wire[35:0] T43;
  wire[17:0] T44;
  reg [17:0] R45;
  reg [17:0] R46;
  wire[17:0] T47;
  reg [17:0] R48;
  reg [17:0] R49;
  wire[17:0] T50;
  wire[17:0] T51;
  wire[17:0] T1138;
  wire[21:0] T52;
  wire[35:0] T53;
  wire[17:0] T54;
  reg [17:0] R55;
  reg [17:0] R56;
  wire[17:0] T57;
  reg [17:0] R58;
  reg [17:0] R59;
  wire T60;
  wire[17:0] T61;
  wire[17:0] T62;
  wire T63;
  wire[17:0] T64;
  wire[17:0] T65;
  wire[17:0] T66;
  wire[17:0] T67;
  wire[17:0] T68;
  wire[17:0] T69;
  wire[17:0] T70;
  wire[17:0] T1139;
  wire[21:0] T71;
  wire[35:0] T72;
  wire[17:0] T73;
  reg [17:0] R74;
  wire[17:0] T75;
  reg [17:0] R76;
  wire[17:0] T77;
  wire[17:0] T78;
  wire[17:0] T79;
  wire[17:0] T80;
  wire[17:0] T81;
  wire[17:0] T1140;
  wire[21:0] T82;
  wire[35:0] T83;
  wire[17:0] T84;
  reg [17:0] R85;
  wire[17:0] T86;
  reg [17:0] R87;
  wire[17:0] T88;
  wire[17:0] T89;
  wire[17:0] T1141;
  wire[21:0] T90;
  wire[35:0] T91;
  wire[17:0] T92;
  reg [17:0] R93;
  wire[17:0] T94;
  reg [17:0] R95;
  wire[17:0] T96;
  reg [17:0] R97;
  reg [17:0] R98;
  wire[17:0] zout_1;
  wire[17:0] T99;
  wire[17:0] T100;
  reg [17:0] R101;
  wire[17:0] T102;
  wire[17:0] T1142;
  wire[21:0] T103;
  wire[35:0] T104;
  wire[17:0] T105;
  wire[17:0] T106;
  wire[17:0] T107;
  wire[17:0] T1143;
  wire[21:0] T108;
  wire[35:0] T109;
  wire[17:0] T110;
  wire[17:0] T111;
  wire[17:0] T112;
  wire[17:0] T113;
  wire[17:0] T114;
  reg [17:0] R115;
  wire[17:0] T116;
  wire[17:0] T117;
  wire[17:0] T118;
  wire[17:0] T119;
  wire[17:0] T120;
  reg [17:0] R121;
  reg [17:0] R122;
  wire[17:0] T123;
  wire[17:0] T124;
  wire[17:0] T125;
  wire[17:0] T126;
  wire[17:0] T127;
  wire[17:0] T1144;
  wire[21:0] T128;
  wire[35:0] T129;
  wire[17:0] T130;
  wire[17:0] T131;
  reg [17:0] R132;
  reg [17:0] R133;
  wire[17:0] T134;
  wire[17:0] T135;
  wire[17:0] T136;
  wire[17:0] T137;
  wire[17:0] T138;
  wire[17:0] T1145;
  wire[21:0] T139;
  wire[35:0] T140;
  wire[17:0] T141;
  wire[17:0] T142;
  reg [17:0] R143;
  reg [17:0] R144;
  wire[17:0] T145;
  wire[17:0] T146;
  wire[17:0] T1146;
  wire[21:0] T147;
  wire[35:0] T148;
  wire[17:0] T149;
  wire[17:0] T150;
  reg [17:0] R151;
  reg [17:0] R152;
  wire T153;
  wire[17:0] T154;
  wire[17:0] T155;
  wire T156;
  wire[17:0] T157;
  wire[17:0] T158;
  wire[17:0] T159;
  wire[17:0] T160;
  wire[17:0] T161;
  wire[17:0] T162;
  wire[17:0] T163;
  wire[17:0] T1147;
  wire[21:0] T164;
  wire[35:0] T165;
  wire[17:0] T166;
  wire[17:0] T167;
  reg [17:0] R168;
  wire[17:0] T169;
  wire[17:0] T170;
  wire[17:0] T171;
  wire[17:0] T172;
  wire[17:0] T173;
  wire[17:0] T1148;
  wire[21:0] T174;
  wire[35:0] T175;
  wire[17:0] T176;
  wire[17:0] T177;
  reg [17:0] R178;
  wire[17:0] T179;
  wire[17:0] T180;
  wire[17:0] T1149;
  wire[21:0] T181;
  wire[35:0] T182;
  wire[17:0] T183;
  wire[17:0] T184;
  reg [17:0] R185;
  wire[17:0] T186;
  reg [17:0] R187;
  reg [17:0] R188;
  wire[17:0] zout_2;
  wire[17:0] T189;
  wire[17:0] T190;
  reg [17:0] R191;
  wire[17:0] T192;
  wire[17:0] T1150;
  wire[21:0] T193;
  wire[35:0] T194;
  wire[17:0] T195;
  wire[17:0] T196;
  wire[17:0] T197;
  wire[17:0] T1151;
  wire[21:0] T198;
  wire[35:0] T199;
  wire[17:0] T200;
  wire[17:0] T201;
  wire[17:0] T202;
  wire[17:0] T203;
  wire[17:0] T204;
  reg [17:0] R205;
  wire[17:0] T206;
  wire[17:0] T207;
  wire[17:0] T208;
  wire[17:0] T209;
  wire[17:0] T210;
  reg [17:0] R211;
  reg [17:0] R212;
  wire[17:0] T213;
  wire[17:0] T214;
  wire[17:0] T215;
  wire[17:0] T216;
  wire[17:0] T217;
  wire[17:0] T1152;
  wire[21:0] T218;
  wire[35:0] T219;
  wire[17:0] T220;
  wire[17:0] T221;
  reg [17:0] R222;
  reg [17:0] R223;
  wire[17:0] T224;
  wire[17:0] T225;
  wire[17:0] T226;
  wire[17:0] T227;
  wire[17:0] T228;
  wire[17:0] T1153;
  wire[21:0] T229;
  wire[35:0] T230;
  wire[17:0] T231;
  wire[17:0] T232;
  reg [17:0] R233;
  reg [17:0] R234;
  wire[17:0] T235;
  wire[17:0] T236;
  wire[17:0] T1154;
  wire[21:0] T237;
  wire[35:0] T238;
  wire[17:0] T239;
  wire[17:0] T240;
  reg [17:0] R241;
  reg [17:0] R242;
  wire T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire T246;
  wire[17:0] T247;
  wire[17:0] T248;
  wire[17:0] T249;
  wire[17:0] T250;
  wire[17:0] T251;
  wire[17:0] T252;
  wire[17:0] T253;
  wire[17:0] T1155;
  wire[21:0] T254;
  wire[35:0] T255;
  wire[17:0] T256;
  wire[17:0] T257;
  reg [17:0] R258;
  wire[17:0] T259;
  wire[17:0] T260;
  wire[17:0] T261;
  wire[17:0] T262;
  wire[17:0] T263;
  wire[17:0] T1156;
  wire[21:0] T264;
  wire[35:0] T265;
  wire[17:0] T266;
  wire[17:0] T267;
  reg [17:0] R268;
  wire[17:0] T269;
  wire[17:0] T270;
  wire[17:0] T1157;
  wire[21:0] T271;
  wire[35:0] T272;
  wire[17:0] T273;
  wire[17:0] T274;
  reg [17:0] R275;
  wire[17:0] T276;
  reg [17:0] R277;
  reg [17:0] R278;
  wire[17:0] yout_0;
  wire[17:0] T279;
  wire[17:0] T280;
  reg [17:0] R281;
  wire[17:0] T282;
  wire[17:0] T1158;
  wire[21:0] T283;
  wire[35:0] T284;
  wire[17:0] T285;
  wire[17:0] T286;
  wire[17:0] T287;
  wire[17:0] T1159;
  wire[21:0] T288;
  wire[35:0] T289;
  wire[17:0] T290;
  wire[17:0] T291;
  wire[17:0] T292;
  wire[17:0] T293;
  wire[17:0] T294;
  reg [17:0] R295;
  reg [17:0] R296;
  reg [17:0] R297;
  wire[17:0] T298;
  reg [17:0] R299;
  reg [17:0] R300;
  wire[17:0] T301;
  wire[17:0] T302;
  wire[17:0] T303;
  wire[17:0] T304;
  wire[17:0] T305;
  wire[17:0] T306;
  wire[17:0] T307;
  wire[17:0] T308;
  wire[17:0] T309;
  reg [17:0] R310;
  wire[17:0] T311;
  wire[17:0] T312;
  wire[17:0] T313;
  wire[17:0] T314;
  wire[17:0] T315;
  wire[17:0] T1160;
  wire[21:0] T316;
  wire[35:0] T317;
  wire[17:0] T318;
  wire[17:0] T319;
  reg [17:0] R320;
  wire[17:0] T321;
  wire[17:0] T322;
  wire[17:0] T323;
  wire[17:0] T324;
  wire[17:0] T325;
  wire[17:0] T1161;
  wire[21:0] T326;
  wire[35:0] T327;
  wire[17:0] T328;
  wire[17:0] T329;
  reg [17:0] R330;
  wire[17:0] T331;
  wire[17:0] T332;
  wire[17:0] T1162;
  wire[21:0] T333;
  wire[35:0] T334;
  wire[17:0] T335;
  wire[17:0] T336;
  reg [17:0] R337;
  wire T338;
  wire[17:0] T339;
  wire[17:0] T340;
  wire T341;
  wire[17:0] T342;
  wire[17:0] T343;
  wire[17:0] T344;
  reg [17:0] R345;
  wire[17:0] yout_1;
  wire[17:0] T346;
  wire[17:0] T347;
  reg [17:0] R348;
  wire[17:0] T349;
  wire[17:0] T1163;
  wire[21:0] T350;
  wire[35:0] T351;
  wire[17:0] T352;
  wire[17:0] T353;
  wire[17:0] T354;
  wire[17:0] T1164;
  wire[21:0] T355;
  wire[35:0] T356;
  wire[17:0] T357;
  wire[17:0] T358;
  wire[17:0] T359;
  wire[17:0] T360;
  wire[17:0] T361;
  reg [17:0] R362;
  reg [17:0] R363;
  reg [17:0] R364;
  wire[17:0] T365;
  reg [17:0] R366;
  reg [17:0] R367;
  wire[17:0] T368;
  wire[17:0] T369;
  wire[17:0] T370;
  wire[17:0] T371;
  wire[17:0] T372;
  wire[17:0] T373;
  wire[17:0] T374;
  wire[17:0] T375;
  wire[17:0] T376;
  reg [17:0] R377;
  wire[17:0] T378;
  wire[17:0] T379;
  wire[17:0] T380;
  wire[17:0] T381;
  wire[17:0] T382;
  wire[17:0] T1165;
  wire[21:0] T383;
  wire[35:0] T384;
  wire[17:0] T385;
  wire[17:0] T386;
  reg [17:0] R387;
  wire[17:0] T388;
  wire[17:0] T389;
  wire[17:0] T390;
  wire[17:0] T391;
  wire[17:0] T392;
  wire[17:0] T1166;
  wire[21:0] T393;
  wire[35:0] T394;
  wire[17:0] T395;
  wire[17:0] T396;
  reg [17:0] R397;
  wire[17:0] T398;
  wire[17:0] T399;
  wire[17:0] T1167;
  wire[21:0] T400;
  wire[35:0] T401;
  wire[17:0] T402;
  wire[17:0] T403;
  reg [17:0] R404;
  wire T405;
  wire[17:0] T406;
  wire[17:0] T407;
  wire T408;
  wire[17:0] T409;
  wire[17:0] T410;
  wire[17:0] T411;
  reg [17:0] R412;
  wire[17:0] yout_2;
  wire[17:0] T413;
  wire[17:0] T414;
  reg [17:0] R415;
  wire[17:0] T416;
  wire[17:0] T1168;
  wire[21:0] T417;
  wire[35:0] T418;
  wire[17:0] T419;
  wire[17:0] T420;
  wire[17:0] T421;
  wire[17:0] T1169;
  wire[21:0] T422;
  wire[35:0] T423;
  wire[17:0] T424;
  wire[17:0] T425;
  wire[17:0] T426;
  wire[17:0] T427;
  wire[17:0] T428;
  reg [17:0] R429;
  reg [17:0] R430;
  reg [17:0] R431;
  wire[17:0] T432;
  reg [17:0] R433;
  reg [17:0] R434;
  wire[17:0] T435;
  wire[17:0] T436;
  wire[17:0] T437;
  wire[17:0] T438;
  wire[17:0] T439;
  wire[17:0] T440;
  wire[17:0] T441;
  wire[17:0] T442;
  wire[17:0] T443;
  reg [17:0] R444;
  wire[17:0] T445;
  wire[17:0] T446;
  wire[17:0] T447;
  wire[17:0] T448;
  wire[17:0] T449;
  wire[17:0] T1170;
  wire[21:0] T450;
  wire[35:0] T451;
  wire[17:0] T452;
  wire[17:0] T453;
  reg [17:0] R454;
  wire[17:0] T455;
  wire[17:0] T456;
  wire[17:0] T457;
  wire[17:0] T458;
  wire[17:0] T459;
  wire[17:0] T1171;
  wire[21:0] T460;
  wire[35:0] T461;
  wire[17:0] T462;
  wire[17:0] T463;
  reg [17:0] R464;
  wire[17:0] T465;
  wire[17:0] T466;
  wire[17:0] T1172;
  wire[21:0] T467;
  wire[35:0] T468;
  wire[17:0] T469;
  wire[17:0] T470;
  reg [17:0] R471;
  wire T472;
  wire[17:0] T473;
  wire[17:0] T474;
  wire T475;
  wire[17:0] T476;
  wire[17:0] T477;
  wire[17:0] T478;
  reg [17:0] R479;
  wire[17:0] yout_3;
  wire[17:0] T480;
  wire[17:0] T481;
  reg [17:0] R482;
  wire[17:0] T483;
  wire[17:0] T1173;
  wire[21:0] T484;
  wire[35:0] T485;
  wire[17:0] T486;
  wire[17:0] T487;
  wire[17:0] T488;
  wire[17:0] T1174;
  wire[21:0] T489;
  wire[35:0] T490;
  wire[17:0] T491;
  wire[17:0] T492;
  wire[17:0] T493;
  wire[17:0] T494;
  wire[17:0] T495;
  reg [17:0] R496;
  reg [17:0] R497;
  reg [17:0] R498;
  wire[17:0] T499;
  reg [17:0] R500;
  reg [17:0] R501;
  wire[17:0] T502;
  wire[17:0] T503;
  wire[17:0] T504;
  wire[17:0] T505;
  wire[17:0] T506;
  wire[17:0] T507;
  wire[17:0] T508;
  wire[17:0] T509;
  wire[17:0] T510;
  reg [17:0] R511;
  wire[17:0] T512;
  wire[17:0] T513;
  wire[17:0] T514;
  wire[17:0] T515;
  wire[17:0] T516;
  wire[17:0] T1175;
  wire[21:0] T517;
  wire[35:0] T518;
  wire[17:0] T519;
  wire[17:0] T520;
  reg [17:0] R521;
  wire[17:0] T522;
  wire[17:0] T523;
  wire[17:0] T524;
  wire[17:0] T525;
  wire[17:0] T526;
  wire[17:0] T1176;
  wire[21:0] T527;
  wire[35:0] T528;
  wire[17:0] T529;
  wire[17:0] T530;
  reg [17:0] R531;
  wire[17:0] T532;
  wire[17:0] T533;
  wire[17:0] T1177;
  wire[21:0] T534;
  wire[35:0] T535;
  wire[17:0] T536;
  wire[17:0] T537;
  reg [17:0] R538;
  wire T539;
  wire[17:0] T540;
  wire[17:0] T541;
  wire T542;
  wire[17:0] T543;
  wire[17:0] T544;
  wire[17:0] T545;
  reg [17:0] R546;
  wire[17:0] yout_4;
  wire[17:0] T547;
  wire[17:0] T548;
  reg [17:0] R549;
  wire[17:0] T550;
  wire[17:0] T1178;
  wire[21:0] T551;
  wire[35:0] T552;
  wire[17:0] T553;
  wire[17:0] T554;
  wire[17:0] T555;
  wire[17:0] T1179;
  wire[21:0] T556;
  wire[35:0] T557;
  wire[17:0] T558;
  wire[17:0] T559;
  wire[17:0] T560;
  wire[17:0] T561;
  wire[17:0] T562;
  reg [17:0] R563;
  reg [17:0] R564;
  reg [17:0] R565;
  wire[17:0] T566;
  reg [17:0] R567;
  reg [17:0] R568;
  wire[17:0] T569;
  wire[17:0] T570;
  wire[17:0] T571;
  wire[17:0] T572;
  wire[17:0] T573;
  wire[17:0] T574;
  wire[17:0] T575;
  wire[17:0] T576;
  wire[17:0] T577;
  reg [17:0] R578;
  wire[17:0] T579;
  wire[17:0] T580;
  wire[17:0] T581;
  wire[17:0] T582;
  wire[17:0] T583;
  wire[17:0] T1180;
  wire[21:0] T584;
  wire[35:0] T585;
  wire[17:0] T586;
  wire[17:0] T587;
  reg [17:0] R588;
  wire[17:0] T589;
  wire[17:0] T590;
  wire[17:0] T591;
  wire[17:0] T592;
  wire[17:0] T593;
  wire[17:0] T1181;
  wire[21:0] T594;
  wire[35:0] T595;
  wire[17:0] T596;
  wire[17:0] T597;
  reg [17:0] R598;
  wire[17:0] T599;
  wire[17:0] T600;
  wire[17:0] T1182;
  wire[21:0] T601;
  wire[35:0] T602;
  wire[17:0] T603;
  wire[17:0] T604;
  reg [17:0] R605;
  wire T606;
  wire[17:0] T607;
  wire[17:0] T608;
  wire T609;
  wire[17:0] T610;
  wire[17:0] T611;
  wire[17:0] T612;
  reg [17:0] R613;
  wire[17:0] yout_5;
  wire[17:0] T614;
  wire[17:0] T615;
  reg [17:0] R616;
  wire[17:0] T617;
  wire[17:0] T1183;
  wire[21:0] T618;
  wire[35:0] T619;
  wire[17:0] T620;
  wire[17:0] T621;
  wire[17:0] T622;
  wire[17:0] T1184;
  wire[21:0] T623;
  wire[35:0] T624;
  wire[17:0] T625;
  wire[17:0] T626;
  wire[17:0] T627;
  wire[17:0] T628;
  wire[17:0] T629;
  reg [17:0] R630;
  reg [17:0] R631;
  reg [17:0] R632;
  wire[17:0] T633;
  reg [17:0] R634;
  reg [17:0] R635;
  wire[17:0] T636;
  wire[17:0] T637;
  wire[17:0] T638;
  wire[17:0] T639;
  wire[17:0] T640;
  wire[17:0] T641;
  wire[17:0] T642;
  wire[17:0] T643;
  wire[17:0] T644;
  reg [17:0] R645;
  wire[17:0] T646;
  wire[17:0] T647;
  wire[17:0] T648;
  wire[17:0] T649;
  wire[17:0] T650;
  wire[17:0] T1185;
  wire[21:0] T651;
  wire[35:0] T652;
  wire[17:0] T653;
  wire[17:0] T654;
  reg [17:0] R655;
  wire[17:0] T656;
  wire[17:0] T657;
  wire[17:0] T658;
  wire[17:0] T659;
  wire[17:0] T660;
  wire[17:0] T1186;
  wire[21:0] T661;
  wire[35:0] T662;
  wire[17:0] T663;
  wire[17:0] T664;
  reg [17:0] R665;
  wire[17:0] T666;
  wire[17:0] T667;
  wire[17:0] T1187;
  wire[21:0] T668;
  wire[35:0] T669;
  wire[17:0] T670;
  wire[17:0] T671;
  reg [17:0] R672;
  wire T673;
  wire[17:0] T674;
  wire[17:0] T675;
  wire T676;
  wire[17:0] T677;
  wire[17:0] T678;
  wire[17:0] T679;
  reg [17:0] R680;
  wire[17:0] yout_6;
  wire[17:0] T681;
  wire[17:0] T682;
  reg [17:0] R683;
  wire[17:0] T684;
  wire[17:0] T1188;
  wire[21:0] T685;
  wire[35:0] T686;
  wire[17:0] T687;
  wire[17:0] T688;
  wire[17:0] T689;
  wire[17:0] T1189;
  wire[21:0] T690;
  wire[35:0] T691;
  wire[17:0] T692;
  wire[17:0] T693;
  wire[17:0] T694;
  wire[17:0] T695;
  wire[17:0] T696;
  reg [17:0] R697;
  reg [17:0] R698;
  reg [17:0] R699;
  wire[17:0] T700;
  reg [17:0] R701;
  reg [17:0] R702;
  wire[17:0] T703;
  wire[17:0] T704;
  wire[17:0] T705;
  wire[17:0] T706;
  wire[17:0] T707;
  wire[17:0] T708;
  wire[17:0] T709;
  wire[17:0] T710;
  wire[17:0] T711;
  reg [17:0] R712;
  wire[17:0] T713;
  wire[17:0] T714;
  wire[17:0] T715;
  wire[17:0] T716;
  wire[17:0] T717;
  wire[17:0] T1190;
  wire[21:0] T718;
  wire[35:0] T719;
  wire[17:0] T720;
  wire[17:0] T721;
  reg [17:0] R722;
  wire[17:0] T723;
  wire[17:0] T724;
  wire[17:0] T725;
  wire[17:0] T726;
  wire[17:0] T727;
  wire[17:0] T1191;
  wire[21:0] T728;
  wire[35:0] T729;
  wire[17:0] T730;
  wire[17:0] T731;
  reg [17:0] R732;
  wire[17:0] T733;
  wire[17:0] T734;
  wire[17:0] T1192;
  wire[21:0] T735;
  wire[35:0] T736;
  wire[17:0] T737;
  wire[17:0] T738;
  reg [17:0] R739;
  wire T740;
  wire[17:0] T741;
  wire[17:0] T742;
  wire T743;
  wire[17:0] T744;
  wire[17:0] T745;
  wire[17:0] T746;
  reg [17:0] R747;
  wire[17:0] yout_7;
  wire[17:0] T748;
  wire[17:0] T749;
  reg [17:0] R750;
  wire[17:0] T751;
  wire[17:0] T1193;
  wire[21:0] T752;
  wire[35:0] T753;
  wire[17:0] T754;
  wire[17:0] T755;
  wire[17:0] T756;
  wire[17:0] T1194;
  wire[21:0] T757;
  wire[35:0] T758;
  wire[17:0] T759;
  wire[17:0] T760;
  wire[17:0] T761;
  wire[17:0] T762;
  wire[17:0] T763;
  reg [17:0] R764;
  reg [17:0] R765;
  reg [17:0] R766;
  wire[17:0] T767;
  reg [17:0] R768;
  reg [17:0] R769;
  wire[17:0] T770;
  wire[17:0] T771;
  wire[17:0] T772;
  wire[17:0] T773;
  wire[17:0] T774;
  wire[17:0] T775;
  wire[17:0] T776;
  wire[17:0] T777;
  wire[17:0] T778;
  reg [17:0] R779;
  wire[17:0] T780;
  wire[17:0] T781;
  wire[17:0] T782;
  wire[17:0] T783;
  wire[17:0] T784;
  wire[17:0] T1195;
  wire[21:0] T785;
  wire[35:0] T786;
  wire[17:0] T787;
  wire[17:0] T788;
  reg [17:0] R789;
  wire[17:0] T790;
  wire[17:0] T791;
  wire[17:0] T792;
  wire[17:0] T793;
  wire[17:0] T794;
  wire[17:0] T1196;
  wire[21:0] T795;
  wire[35:0] T796;
  wire[17:0] T797;
  wire[17:0] T798;
  reg [17:0] R799;
  wire[17:0] T800;
  wire[17:0] T801;
  wire[17:0] T1197;
  wire[21:0] T802;
  wire[35:0] T803;
  wire[17:0] T804;
  wire[17:0] T805;
  reg [17:0] R806;
  wire T807;
  wire[17:0] T808;
  wire[17:0] T809;
  wire T810;
  wire[17:0] T811;
  wire[17:0] T812;
  wire[17:0] T813;
  reg [17:0] R814;
  wire[17:0] yout_8;
  wire[17:0] T815;
  wire[17:0] T816;
  reg [17:0] R817;
  wire[17:0] T818;
  wire[17:0] T1198;
  wire[21:0] T819;
  wire[35:0] T820;
  wire[17:0] T821;
  wire[17:0] T822;
  wire[17:0] T823;
  wire[17:0] T1199;
  wire[21:0] T824;
  wire[35:0] T825;
  wire[17:0] T826;
  wire[17:0] T827;
  wire[17:0] T828;
  wire[17:0] T829;
  wire[17:0] T830;
  reg [17:0] R831;
  reg [17:0] R832;
  reg [17:0] R833;
  wire[17:0] T834;
  reg [17:0] R835;
  reg [17:0] R836;
  wire[17:0] T837;
  wire[17:0] T838;
  wire[17:0] T839;
  wire[17:0] T840;
  wire[17:0] T841;
  wire[17:0] T842;
  wire[17:0] T843;
  wire[17:0] T844;
  wire[17:0] T845;
  reg [17:0] R846;
  wire[17:0] T847;
  wire[17:0] T848;
  wire[17:0] T849;
  wire[17:0] T850;
  wire[17:0] T851;
  wire[17:0] T1200;
  wire[21:0] T852;
  wire[35:0] T853;
  wire[17:0] T854;
  wire[17:0] T855;
  reg [17:0] R856;
  wire[17:0] T857;
  wire[17:0] T858;
  wire[17:0] T859;
  wire[17:0] T860;
  wire[17:0] T861;
  wire[17:0] T1201;
  wire[21:0] T862;
  wire[35:0] T863;
  wire[17:0] T864;
  wire[17:0] T865;
  reg [17:0] R866;
  wire[17:0] T867;
  wire[17:0] T868;
  wire[17:0] T1202;
  wire[21:0] T869;
  wire[35:0] T870;
  wire[17:0] T871;
  wire[17:0] T872;
  reg [17:0] R873;
  wire T874;
  wire[17:0] T875;
  wire[17:0] T876;
  wire T877;
  wire[17:0] T878;
  wire[17:0] T879;
  wire[17:0] T880;
  reg [17:0] R881;
  wire[17:0] yout_9;
  wire[17:0] T882;
  wire[17:0] T883;
  reg [17:0] R884;
  wire[17:0] T885;
  wire[17:0] T1203;
  wire[21:0] T886;
  wire[35:0] T887;
  wire[17:0] T888;
  wire[17:0] T889;
  wire[17:0] T890;
  wire[17:0] T1204;
  wire[21:0] T891;
  wire[35:0] T892;
  wire[17:0] T893;
  wire[17:0] T894;
  wire[17:0] T895;
  wire[17:0] T896;
  wire[17:0] T897;
  reg [17:0] R898;
  reg [17:0] R899;
  reg [17:0] R900;
  wire[17:0] T901;
  reg [17:0] R902;
  reg [17:0] R903;
  wire[17:0] T904;
  wire[17:0] T905;
  wire[17:0] T906;
  wire[17:0] T907;
  wire[17:0] T908;
  wire[17:0] T909;
  wire[17:0] T910;
  wire[17:0] T911;
  wire[17:0] T912;
  reg [17:0] R913;
  wire[17:0] T914;
  wire[17:0] T915;
  wire[17:0] T916;
  wire[17:0] T917;
  wire[17:0] T918;
  wire[17:0] T1205;
  wire[21:0] T919;
  wire[35:0] T920;
  wire[17:0] T921;
  wire[17:0] T922;
  reg [17:0] R923;
  wire[17:0] T924;
  wire[17:0] T925;
  wire[17:0] T926;
  wire[17:0] T927;
  wire[17:0] T928;
  wire[17:0] T1206;
  wire[21:0] T929;
  wire[35:0] T930;
  wire[17:0] T931;
  wire[17:0] T932;
  reg [17:0] R933;
  wire[17:0] T934;
  wire[17:0] T935;
  wire[17:0] T1207;
  wire[21:0] T936;
  wire[35:0] T937;
  wire[17:0] T938;
  wire[17:0] T939;
  reg [17:0] R940;
  wire T941;
  wire[17:0] T942;
  wire[17:0] T943;
  wire T944;
  wire[17:0] T945;
  wire[17:0] T946;
  wire[17:0] T947;
  reg [17:0] R948;
  wire[17:0] yout_10;
  wire[17:0] T949;
  wire[17:0] T950;
  reg [17:0] R951;
  wire[17:0] T952;
  wire[17:0] T1208;
  wire[21:0] T953;
  wire[35:0] T954;
  wire[17:0] T955;
  wire[17:0] T956;
  wire[17:0] T957;
  wire[17:0] T1209;
  wire[21:0] T958;
  wire[35:0] T959;
  wire[17:0] T960;
  wire[17:0] T961;
  wire[17:0] T962;
  wire[17:0] T963;
  wire[17:0] T964;
  reg [17:0] R965;
  reg [17:0] R966;
  reg [17:0] R967;
  wire[17:0] T968;
  reg [17:0] R969;
  reg [17:0] R970;
  wire[17:0] T971;
  wire[17:0] T972;
  wire[17:0] T973;
  wire[17:0] T974;
  wire[17:0] T975;
  wire[17:0] T976;
  wire[17:0] T977;
  wire[17:0] T978;
  wire[17:0] T979;
  reg [17:0] R980;
  wire[17:0] T981;
  wire[17:0] T982;
  wire[17:0] T983;
  wire[17:0] T984;
  wire[17:0] T985;
  wire[17:0] T1210;
  wire[21:0] T986;
  wire[35:0] T987;
  wire[17:0] T988;
  wire[17:0] T989;
  reg [17:0] R990;
  wire[17:0] T991;
  wire[17:0] T992;
  wire[17:0] T993;
  wire[17:0] T994;
  wire[17:0] T995;
  wire[17:0] T1211;
  wire[21:0] T996;
  wire[35:0] T997;
  wire[17:0] T998;
  wire[17:0] T999;
  reg [17:0] R1000;
  wire[17:0] T1001;
  wire[17:0] T1002;
  wire[17:0] T1212;
  wire[21:0] T1003;
  wire[35:0] T1004;
  wire[17:0] T1005;
  wire[17:0] T1006;
  reg [17:0] R1007;
  wire T1008;
  wire[17:0] T1009;
  wire[17:0] T1010;
  wire T1011;
  wire[17:0] T1012;
  wire[17:0] T1013;
  wire[17:0] T1014;
  reg [17:0] R1015;
  wire[17:0] yout_11;
  wire[17:0] T1016;
  wire[17:0] T1017;
  reg [17:0] R1018;
  wire[17:0] T1019;
  wire[17:0] T1213;
  wire[21:0] T1020;
  wire[35:0] T1021;
  wire[17:0] T1022;
  wire[17:0] T1023;
  wire[17:0] T1024;
  wire[17:0] T1214;
  wire[21:0] T1025;
  wire[35:0] T1026;
  wire[17:0] T1027;
  wire[17:0] T1028;
  wire[17:0] T1029;
  wire[17:0] T1030;
  wire[17:0] T1031;
  reg [17:0] R1032;
  reg [17:0] R1033;
  reg [17:0] R1034;
  wire[17:0] T1035;
  reg [17:0] R1036;
  reg [17:0] R1037;
  wire[17:0] T1038;
  wire[17:0] T1039;
  wire[17:0] T1040;
  wire[17:0] T1041;
  wire[17:0] T1042;
  wire[17:0] T1043;
  wire[17:0] T1044;
  wire[17:0] T1045;
  wire[17:0] T1046;
  reg [17:0] R1047;
  wire[17:0] T1048;
  wire[17:0] T1049;
  wire[17:0] T1050;
  wire[17:0] T1051;
  wire[17:0] T1052;
  wire[17:0] T1215;
  wire[21:0] T1053;
  wire[35:0] T1054;
  wire[17:0] T1055;
  wire[17:0] T1056;
  reg [17:0] R1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[17:0] T1060;
  wire[17:0] T1061;
  wire[17:0] T1062;
  wire[17:0] T1216;
  wire[21:0] T1063;
  wire[35:0] T1064;
  wire[17:0] T1065;
  wire[17:0] T1066;
  reg [17:0] R1067;
  wire[17:0] T1068;
  wire[17:0] T1069;
  wire[17:0] T1217;
  wire[21:0] T1070;
  wire[35:0] T1071;
  wire[17:0] T1072;
  wire[17:0] T1073;
  reg [17:0] R1074;
  wire T1075;
  wire[17:0] T1076;
  wire[17:0] T1077;
  wire T1078;
  wire[17:0] T1079;
  wire[17:0] T1080;
  wire[17:0] T1081;
  reg [17:0] R1082;
  wire[17:0] xout_0;
  wire[17:0] T1083;
  wire[17:0] T1084;
  reg [17:0] R1085;
  wire[17:0] T1086;
  wire[17:0] T1218;
  wire[21:0] T1087;
  wire[35:0] T1088;
  wire[17:0] T1089;
  wire[17:0] T1090;
  wire[17:0] T1091;
  wire[17:0] T1092;
  wire[17:0] T1093;
  reg [17:0] R1094;
  reg [17:0] R1095;
  reg [17:0] R1096;
  wire[17:0] T1097;
  wire[17:0] T1098;
  reg [17:0] R1099;
  wire[17:0] xout_1;
  wire[17:0] T1100;
  wire[17:0] T1101;
  reg [17:0] R1102;
  wire[17:0] T1103;
  wire[17:0] T1219;
  wire[21:0] T1104;
  wire[35:0] T1105;
  wire[17:0] T1106;
  wire[17:0] T1107;
  wire[17:0] T1108;
  wire[17:0] T1109;
  wire[17:0] T1110;
  reg [17:0] R1111;
  reg [17:0] R1112;
  reg [17:0] R1113;
  wire[17:0] T1114;
  wire[17:0] T1115;
  reg [17:0] R1116;
  wire[17:0] xout_2;
  wire[17:0] T1117;
  wire[17:0] T1118;
  reg [17:0] R1119;
  wire[17:0] T1120;
  wire[17:0] T1220;
  wire[21:0] T1121;
  wire[35:0] T1122;
  wire[17:0] T1123;
  wire[17:0] T1124;
  wire[17:0] T1125;
  wire[17:0] T1126;
  wire[17:0] T1127;
  reg [17:0] R1128;
  reg [17:0] R1129;
  reg [17:0] R1130;
  wire[17:0] T1131;
  wire[17:0] T1132;
  reg [17:0] R1133;
  wire[17:0] XNetModule_io_o_2;
  wire[17:0] XNetModule_io_o_1;
  wire[17:0] XNetModule_io_o_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R2 = {1{$random}};
    R16 = {1{$random}};
    R22 = {1{$random}};
    R23 = {1{$random}};
    R32 = {1{$random}};
    R33 = {1{$random}};
    R35 = {1{$random}};
    R36 = {1{$random}};
    R45 = {1{$random}};
    R46 = {1{$random}};
    R48 = {1{$random}};
    R49 = {1{$random}};
    R55 = {1{$random}};
    R56 = {1{$random}};
    R58 = {1{$random}};
    R59 = {1{$random}};
    R74 = {1{$random}};
    R76 = {1{$random}};
    R85 = {1{$random}};
    R87 = {1{$random}};
    R93 = {1{$random}};
    R95 = {1{$random}};
    R97 = {1{$random}};
    R98 = {1{$random}};
    R101 = {1{$random}};
    R115 = {1{$random}};
    R121 = {1{$random}};
    R122 = {1{$random}};
    R132 = {1{$random}};
    R133 = {1{$random}};
    R143 = {1{$random}};
    R144 = {1{$random}};
    R151 = {1{$random}};
    R152 = {1{$random}};
    R168 = {1{$random}};
    R178 = {1{$random}};
    R185 = {1{$random}};
    R187 = {1{$random}};
    R188 = {1{$random}};
    R191 = {1{$random}};
    R205 = {1{$random}};
    R211 = {1{$random}};
    R212 = {1{$random}};
    R222 = {1{$random}};
    R223 = {1{$random}};
    R233 = {1{$random}};
    R234 = {1{$random}};
    R241 = {1{$random}};
    R242 = {1{$random}};
    R258 = {1{$random}};
    R268 = {1{$random}};
    R275 = {1{$random}};
    R277 = {1{$random}};
    R278 = {1{$random}};
    R281 = {1{$random}};
    R295 = {1{$random}};
    R296 = {1{$random}};
    R297 = {1{$random}};
    R299 = {1{$random}};
    R300 = {1{$random}};
    R310 = {1{$random}};
    R320 = {1{$random}};
    R330 = {1{$random}};
    R337 = {1{$random}};
    R345 = {1{$random}};
    R348 = {1{$random}};
    R362 = {1{$random}};
    R363 = {1{$random}};
    R364 = {1{$random}};
    R366 = {1{$random}};
    R367 = {1{$random}};
    R377 = {1{$random}};
    R387 = {1{$random}};
    R397 = {1{$random}};
    R404 = {1{$random}};
    R412 = {1{$random}};
    R415 = {1{$random}};
    R429 = {1{$random}};
    R430 = {1{$random}};
    R431 = {1{$random}};
    R433 = {1{$random}};
    R434 = {1{$random}};
    R444 = {1{$random}};
    R454 = {1{$random}};
    R464 = {1{$random}};
    R471 = {1{$random}};
    R479 = {1{$random}};
    R482 = {1{$random}};
    R496 = {1{$random}};
    R497 = {1{$random}};
    R498 = {1{$random}};
    R500 = {1{$random}};
    R501 = {1{$random}};
    R511 = {1{$random}};
    R521 = {1{$random}};
    R531 = {1{$random}};
    R538 = {1{$random}};
    R546 = {1{$random}};
    R549 = {1{$random}};
    R563 = {1{$random}};
    R564 = {1{$random}};
    R565 = {1{$random}};
    R567 = {1{$random}};
    R568 = {1{$random}};
    R578 = {1{$random}};
    R588 = {1{$random}};
    R598 = {1{$random}};
    R605 = {1{$random}};
    R613 = {1{$random}};
    R616 = {1{$random}};
    R630 = {1{$random}};
    R631 = {1{$random}};
    R632 = {1{$random}};
    R634 = {1{$random}};
    R635 = {1{$random}};
    R645 = {1{$random}};
    R655 = {1{$random}};
    R665 = {1{$random}};
    R672 = {1{$random}};
    R680 = {1{$random}};
    R683 = {1{$random}};
    R697 = {1{$random}};
    R698 = {1{$random}};
    R699 = {1{$random}};
    R701 = {1{$random}};
    R702 = {1{$random}};
    R712 = {1{$random}};
    R722 = {1{$random}};
    R732 = {1{$random}};
    R739 = {1{$random}};
    R747 = {1{$random}};
    R750 = {1{$random}};
    R764 = {1{$random}};
    R765 = {1{$random}};
    R766 = {1{$random}};
    R768 = {1{$random}};
    R769 = {1{$random}};
    R779 = {1{$random}};
    R789 = {1{$random}};
    R799 = {1{$random}};
    R806 = {1{$random}};
    R814 = {1{$random}};
    R817 = {1{$random}};
    R831 = {1{$random}};
    R832 = {1{$random}};
    R833 = {1{$random}};
    R835 = {1{$random}};
    R836 = {1{$random}};
    R846 = {1{$random}};
    R856 = {1{$random}};
    R866 = {1{$random}};
    R873 = {1{$random}};
    R881 = {1{$random}};
    R884 = {1{$random}};
    R898 = {1{$random}};
    R899 = {1{$random}};
    R900 = {1{$random}};
    R902 = {1{$random}};
    R903 = {1{$random}};
    R913 = {1{$random}};
    R923 = {1{$random}};
    R933 = {1{$random}};
    R940 = {1{$random}};
    R948 = {1{$random}};
    R951 = {1{$random}};
    R965 = {1{$random}};
    R966 = {1{$random}};
    R967 = {1{$random}};
    R969 = {1{$random}};
    R970 = {1{$random}};
    R980 = {1{$random}};
    R990 = {1{$random}};
    R1000 = {1{$random}};
    R1007 = {1{$random}};
    R1015 = {1{$random}};
    R1018 = {1{$random}};
    R1032 = {1{$random}};
    R1033 = {1{$random}};
    R1034 = {1{$random}};
    R1036 = {1{$random}};
    R1037 = {1{$random}};
    R1047 = {1{$random}};
    R1057 = {1{$random}};
    R1067 = {1{$random}};
    R1074 = {1{$random}};
    R1082 = {1{$random}};
    R1085 = {1{$random}};
    R1094 = {1{$random}};
    R1095 = {1{$random}};
    R1096 = {1{$random}};
    R1099 = {1{$random}};
    R1102 = {1{$random}};
    R1111 = {1{$random}};
    R1112 = {1{$random}};
    R1113 = {1{$random}};
    R1116 = {1{$random}};
    R1119 = {1{$random}};
    R1128 = {1{$random}};
    R1129 = {1{$random}};
    R1130 = {1{$random}};
    R1133 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_zout_0 = zout_0;
  assign zout_0 = T0;
  assign T0 = T96 + T1;
  assign T1 = R2;
  assign T3 = T1134;
  assign T1134 = T4[5'h11:1'h0];
  assign T4 = $signed(T5) >>> 4'he;
  assign T5 = $signed(T7) * $signed(T6);
  assign T6 = 18'h8000;
  assign T7 = T8;
  assign T8 = T1135;
  assign T1135 = T9[5'h11:1'h0];
  assign T9 = $signed(T10) >>> 4'he;
  assign T10 = $signed(T12) * $signed(T11);
  assign T11 = io_lbda;
  assign T12 = T13;
  assign T13 = T14;
  assign T14 = T66 - T15;
  assign T15 = R16;
  assign T17 = T63 ? 18'h8000 : T18;
  assign T18 = T60 ? 18'h38000 : T19;
  assign T19 = T20;
  assign T20 = T24 - T21;
  assign T21 = R22;
  assign T24 = T25;
  assign T25 = T26;
  assign T26 = T37 + T27;
  assign T27 = T28;
  assign T28 = T1136;
  assign T1136 = T29[5'h11:1'h0];
  assign T29 = $signed(T30) >>> 4'he;
  assign T30 = $signed(T34) * $signed(T31);
  assign T31 = R32;
  assign T34 = R35;
  assign T37 = T38;
  assign T38 = T39;
  assign T39 = T50 + T40;
  assign T40 = T41;
  assign T41 = T1137;
  assign T1137 = T42[5'h11:1'h0];
  assign T42 = $signed(T43) >>> 4'he;
  assign T43 = $signed(T47) * $signed(T44);
  assign T44 = R45;
  assign T47 = R48;
  assign T50 = T51;
  assign T51 = T1138;
  assign T1138 = T52[5'h11:1'h0];
  assign T52 = $signed(T53) >>> 4'he;
  assign T53 = $signed(T57) * $signed(T54);
  assign T54 = R55;
  assign T57 = R58;
  assign T60 = $signed(T62) < $signed(T61);
  assign T61 = 18'h38000;
  assign T62 = T19;
  assign T63 = $signed(T65) < $signed(T64);
  assign T64 = T19;
  assign T65 = 18'h8000;
  assign T66 = T67;
  assign T67 = T68;
  assign T68 = T77 + T69;
  assign T69 = T70;
  assign T70 = T1139;
  assign T1139 = T71[5'h11:1'h0];
  assign T71 = $signed(T72) >>> 4'he;
  assign T72 = $signed(T75) * $signed(T73);
  assign T73 = R74;
  assign T75 = R76;
  assign T77 = T78;
  assign T78 = T79;
  assign T79 = T88 + T80;
  assign T80 = T81;
  assign T81 = T1140;
  assign T1140 = T82[5'h11:1'h0];
  assign T82 = $signed(T83) >>> 4'he;
  assign T83 = $signed(T86) * $signed(T84);
  assign T84 = R85;
  assign T86 = R87;
  assign T88 = T89;
  assign T89 = T1141;
  assign T1141 = T90[5'h11:1'h0];
  assign T90 = $signed(T91) >>> 4'he;
  assign T91 = $signed(T94) * $signed(T92);
  assign T92 = R93;
  assign T94 = R95;
  assign T96 = R97;
  assign io_zout_1 = zout_1;
  assign zout_1 = T99;
  assign T99 = T186 + T100;
  assign T100 = R101;
  assign T102 = T1142;
  assign T1142 = T103[5'h11:1'h0];
  assign T103 = $signed(T104) >>> 4'he;
  assign T104 = $signed(T106) * $signed(T105);
  assign T105 = 18'h8000;
  assign T106 = T107;
  assign T107 = T1143;
  assign T1143 = T108[5'h11:1'h0];
  assign T108 = $signed(T109) >>> 4'he;
  assign T109 = $signed(T111) * $signed(T110);
  assign T110 = io_lbda;
  assign T111 = T112;
  assign T112 = T113;
  assign T113 = T159 - T114;
  assign T114 = R115;
  assign T116 = T156 ? 18'h8000 : T117;
  assign T117 = T153 ? 18'h38000 : T118;
  assign T118 = T119;
  assign T119 = T123 - T120;
  assign T120 = R121;
  assign T123 = T124;
  assign T124 = T125;
  assign T125 = T134 + T126;
  assign T126 = T127;
  assign T127 = T1144;
  assign T1144 = T128[5'h11:1'h0];
  assign T128 = $signed(T129) >>> 4'he;
  assign T129 = $signed(T131) * $signed(T130);
  assign T130 = R32;
  assign T131 = R132;
  assign T134 = T135;
  assign T135 = T136;
  assign T136 = T145 + T137;
  assign T137 = T138;
  assign T138 = T1145;
  assign T1145 = T139[5'h11:1'h0];
  assign T139 = $signed(T140) >>> 4'he;
  assign T140 = $signed(T142) * $signed(T141);
  assign T141 = R45;
  assign T142 = R143;
  assign T145 = T146;
  assign T146 = T1146;
  assign T1146 = T147[5'h11:1'h0];
  assign T147 = $signed(T148) >>> 4'he;
  assign T148 = $signed(T150) * $signed(T149);
  assign T149 = R55;
  assign T150 = R151;
  assign T153 = $signed(T155) < $signed(T154);
  assign T154 = 18'h38000;
  assign T155 = T118;
  assign T156 = $signed(T158) < $signed(T157);
  assign T157 = T118;
  assign T158 = 18'h8000;
  assign T159 = T160;
  assign T160 = T161;
  assign T161 = T169 + T162;
  assign T162 = T163;
  assign T163 = T1147;
  assign T1147 = T164[5'h11:1'h0];
  assign T164 = $signed(T165) >>> 4'he;
  assign T165 = $signed(T167) * $signed(T166);
  assign T166 = R74;
  assign T167 = R168;
  assign T169 = T170;
  assign T170 = T171;
  assign T171 = T179 + T172;
  assign T172 = T173;
  assign T173 = T1148;
  assign T1148 = T174[5'h11:1'h0];
  assign T174 = $signed(T175) >>> 4'he;
  assign T175 = $signed(T177) * $signed(T176);
  assign T176 = R85;
  assign T177 = R178;
  assign T179 = T180;
  assign T180 = T1149;
  assign T1149 = T181[5'h11:1'h0];
  assign T181 = $signed(T182) >>> 4'he;
  assign T182 = $signed(T184) * $signed(T183);
  assign T183 = R93;
  assign T184 = R185;
  assign T186 = R187;
  assign io_zout_2 = zout_2;
  assign zout_2 = T189;
  assign T189 = T276 + T190;
  assign T190 = R191;
  assign T192 = T1150;
  assign T1150 = T193[5'h11:1'h0];
  assign T193 = $signed(T194) >>> 4'he;
  assign T194 = $signed(T196) * $signed(T195);
  assign T195 = 18'h8000;
  assign T196 = T197;
  assign T197 = T1151;
  assign T1151 = T198[5'h11:1'h0];
  assign T198 = $signed(T199) >>> 4'he;
  assign T199 = $signed(T201) * $signed(T200);
  assign T200 = io_lbda;
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = T249 - T204;
  assign T204 = R205;
  assign T206 = T246 ? 18'h8000 : T207;
  assign T207 = T243 ? 18'h38000 : T208;
  assign T208 = T209;
  assign T209 = T213 - T210;
  assign T210 = R211;
  assign T213 = T214;
  assign T214 = T215;
  assign T215 = T224 + T216;
  assign T216 = T217;
  assign T217 = T1152;
  assign T1152 = T218[5'h11:1'h0];
  assign T218 = $signed(T219) >>> 4'he;
  assign T219 = $signed(T221) * $signed(T220);
  assign T220 = R32;
  assign T221 = R222;
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T235 + T227;
  assign T227 = T228;
  assign T228 = T1153;
  assign T1153 = T229[5'h11:1'h0];
  assign T229 = $signed(T230) >>> 4'he;
  assign T230 = $signed(T232) * $signed(T231);
  assign T231 = R45;
  assign T232 = R233;
  assign T235 = T236;
  assign T236 = T1154;
  assign T1154 = T237[5'h11:1'h0];
  assign T237 = $signed(T238) >>> 4'he;
  assign T238 = $signed(T240) * $signed(T239);
  assign T239 = R55;
  assign T240 = R241;
  assign T243 = $signed(T245) < $signed(T244);
  assign T244 = 18'h38000;
  assign T245 = T208;
  assign T246 = $signed(T248) < $signed(T247);
  assign T247 = T208;
  assign T248 = 18'h8000;
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = T259 + T252;
  assign T252 = T253;
  assign T253 = T1155;
  assign T1155 = T254[5'h11:1'h0];
  assign T254 = $signed(T255) >>> 4'he;
  assign T255 = $signed(T257) * $signed(T256);
  assign T256 = R74;
  assign T257 = R258;
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = T269 + T262;
  assign T262 = T263;
  assign T263 = T1156;
  assign T1156 = T264[5'h11:1'h0];
  assign T264 = $signed(T265) >>> 4'he;
  assign T265 = $signed(T267) * $signed(T266);
  assign T266 = R85;
  assign T267 = R268;
  assign T269 = T270;
  assign T270 = T1157;
  assign T1157 = T271[5'h11:1'h0];
  assign T271 = $signed(T272) >>> 4'he;
  assign T272 = $signed(T274) * $signed(T273);
  assign T273 = R93;
  assign T274 = R275;
  assign T276 = R277;
  assign io_yout_0 = yout_0;
  assign yout_0 = T279;
  assign T279 = T344 + T280;
  assign T280 = R281;
  assign T282 = T1158;
  assign T1158 = T283[5'h11:1'h0];
  assign T283 = $signed(T284) >>> 4'he;
  assign T284 = $signed(T286) * $signed(T285);
  assign T285 = 18'h8000;
  assign T286 = T287;
  assign T287 = T1159;
  assign T1159 = T288[5'h11:1'h0];
  assign T288 = $signed(T289) >>> 4'he;
  assign T289 = $signed(T291) * $signed(T290);
  assign T290 = io_lbda;
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = T298 - T294;
  assign T294 = R295;
  assign T298 = R299;
  assign T301 = T341 ? 18'h8000 : T302;
  assign T302 = T338 ? 18'h38000 : T303;
  assign T303 = T304;
  assign T304 = T306 + T305;
  assign T305 = R297;
  assign T306 = T307;
  assign T307 = T308;
  assign T308 = T311 - T309;
  assign T309 = R310;
  assign T311 = T312;
  assign T312 = T313;
  assign T313 = T321 + T314;
  assign T314 = T315;
  assign T315 = T1160;
  assign T1160 = T316[5'h11:1'h0];
  assign T316 = $signed(T317) >>> 4'he;
  assign T317 = $signed(T319) * $signed(T318);
  assign T318 = R33;
  assign T319 = R320;
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = T331 + T324;
  assign T324 = T325;
  assign T325 = T1161;
  assign T1161 = T326[5'h11:1'h0];
  assign T326 = $signed(T327) >>> 4'he;
  assign T327 = $signed(T329) * $signed(T328);
  assign T328 = R46;
  assign T329 = R330;
  assign T331 = T332;
  assign T332 = T1162;
  assign T1162 = T333[5'h11:1'h0];
  assign T333 = $signed(T334) >>> 4'he;
  assign T334 = $signed(T336) * $signed(T335);
  assign T335 = R56;
  assign T336 = R337;
  assign T338 = $signed(T340) < $signed(T339);
  assign T339 = 18'h38000;
  assign T340 = T303;
  assign T341 = $signed(T343) < $signed(T342);
  assign T342 = T303;
  assign T343 = 18'h8000;
  assign T344 = R345;
  assign io_yout_1 = yout_1;
  assign yout_1 = T346;
  assign T346 = T411 + T347;
  assign T347 = R348;
  assign T349 = T1163;
  assign T1163 = T350[5'h11:1'h0];
  assign T350 = $signed(T351) >>> 4'he;
  assign T351 = $signed(T353) * $signed(T352);
  assign T352 = 18'h8000;
  assign T353 = T354;
  assign T354 = T1164;
  assign T1164 = T355[5'h11:1'h0];
  assign T355 = $signed(T356) >>> 4'he;
  assign T356 = $signed(T358) * $signed(T357);
  assign T357 = io_lbda;
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T365 - T361;
  assign T361 = R362;
  assign T365 = R366;
  assign T368 = T408 ? 18'h8000 : T369;
  assign T369 = T405 ? 18'h38000 : T370;
  assign T370 = T371;
  assign T371 = T373 + T372;
  assign T372 = R364;
  assign T373 = T374;
  assign T374 = T375;
  assign T375 = T378 - T376;
  assign T376 = R377;
  assign T378 = T379;
  assign T379 = T380;
  assign T380 = T388 + T381;
  assign T381 = T382;
  assign T382 = T1165;
  assign T1165 = T383[5'h11:1'h0];
  assign T383 = $signed(T384) >>> 4'he;
  assign T384 = $signed(T386) * $signed(T385);
  assign T385 = R33;
  assign T386 = R387;
  assign T388 = T389;
  assign T389 = T390;
  assign T390 = T398 + T391;
  assign T391 = T392;
  assign T392 = T1166;
  assign T1166 = T393[5'h11:1'h0];
  assign T393 = $signed(T394) >>> 4'he;
  assign T394 = $signed(T396) * $signed(T395);
  assign T395 = R46;
  assign T396 = R397;
  assign T398 = T399;
  assign T399 = T1167;
  assign T1167 = T400[5'h11:1'h0];
  assign T400 = $signed(T401) >>> 4'he;
  assign T401 = $signed(T403) * $signed(T402);
  assign T402 = R56;
  assign T403 = R404;
  assign T405 = $signed(T407) < $signed(T406);
  assign T406 = 18'h38000;
  assign T407 = T370;
  assign T408 = $signed(T410) < $signed(T409);
  assign T409 = T370;
  assign T410 = 18'h8000;
  assign T411 = R412;
  assign io_yout_2 = yout_2;
  assign yout_2 = T413;
  assign T413 = T478 + T414;
  assign T414 = R415;
  assign T416 = T1168;
  assign T1168 = T417[5'h11:1'h0];
  assign T417 = $signed(T418) >>> 4'he;
  assign T418 = $signed(T420) * $signed(T419);
  assign T419 = 18'h8000;
  assign T420 = T421;
  assign T421 = T1169;
  assign T1169 = T422[5'h11:1'h0];
  assign T422 = $signed(T423) >>> 4'he;
  assign T423 = $signed(T425) * $signed(T424);
  assign T424 = io_lbda;
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = T432 - T428;
  assign T428 = R429;
  assign T432 = R433;
  assign T435 = T475 ? 18'h8000 : T436;
  assign T436 = T472 ? 18'h38000 : T437;
  assign T437 = T438;
  assign T438 = T440 + T439;
  assign T439 = R431;
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T445 - T443;
  assign T443 = R444;
  assign T445 = T446;
  assign T446 = T447;
  assign T447 = T455 + T448;
  assign T448 = T449;
  assign T449 = T1170;
  assign T1170 = T450[5'h11:1'h0];
  assign T450 = $signed(T451) >>> 4'he;
  assign T451 = $signed(T453) * $signed(T452);
  assign T452 = R33;
  assign T453 = R454;
  assign T455 = T456;
  assign T456 = T457;
  assign T457 = T465 + T458;
  assign T458 = T459;
  assign T459 = T1171;
  assign T1171 = T460[5'h11:1'h0];
  assign T460 = $signed(T461) >>> 4'he;
  assign T461 = $signed(T463) * $signed(T462);
  assign T462 = R46;
  assign T463 = R464;
  assign T465 = T466;
  assign T466 = T1172;
  assign T1172 = T467[5'h11:1'h0];
  assign T467 = $signed(T468) >>> 4'he;
  assign T468 = $signed(T470) * $signed(T469);
  assign T469 = R56;
  assign T470 = R471;
  assign T472 = $signed(T474) < $signed(T473);
  assign T473 = 18'h38000;
  assign T474 = T437;
  assign T475 = $signed(T477) < $signed(T476);
  assign T476 = T437;
  assign T477 = 18'h8000;
  assign T478 = R479;
  assign io_yout_3 = yout_3;
  assign yout_3 = T480;
  assign T480 = T545 + T481;
  assign T481 = R482;
  assign T483 = T1173;
  assign T1173 = T484[5'h11:1'h0];
  assign T484 = $signed(T485) >>> 4'he;
  assign T485 = $signed(T487) * $signed(T486);
  assign T486 = 18'h8000;
  assign T487 = T488;
  assign T488 = T1174;
  assign T1174 = T489[5'h11:1'h0];
  assign T489 = $signed(T490) >>> 4'he;
  assign T490 = $signed(T492) * $signed(T491);
  assign T491 = io_lbda;
  assign T492 = T493;
  assign T493 = T494;
  assign T494 = T499 - T495;
  assign T495 = R496;
  assign T499 = R500;
  assign T502 = T542 ? 18'h8000 : T503;
  assign T503 = T539 ? 18'h38000 : T504;
  assign T504 = T505;
  assign T505 = T507 + T506;
  assign T506 = R498;
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = T512 - T510;
  assign T510 = R511;
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T522 + T515;
  assign T515 = T516;
  assign T516 = T1175;
  assign T1175 = T517[5'h11:1'h0];
  assign T517 = $signed(T518) >>> 4'he;
  assign T518 = $signed(T520) * $signed(T519);
  assign T519 = R33;
  assign T520 = R521;
  assign T522 = T523;
  assign T523 = T524;
  assign T524 = T532 + T525;
  assign T525 = T526;
  assign T526 = T1176;
  assign T1176 = T527[5'h11:1'h0];
  assign T527 = $signed(T528) >>> 4'he;
  assign T528 = $signed(T530) * $signed(T529);
  assign T529 = R46;
  assign T530 = R531;
  assign T532 = T533;
  assign T533 = T1177;
  assign T1177 = T534[5'h11:1'h0];
  assign T534 = $signed(T535) >>> 4'he;
  assign T535 = $signed(T537) * $signed(T536);
  assign T536 = R56;
  assign T537 = R538;
  assign T539 = $signed(T541) < $signed(T540);
  assign T540 = 18'h38000;
  assign T541 = T504;
  assign T542 = $signed(T544) < $signed(T543);
  assign T543 = T504;
  assign T544 = 18'h8000;
  assign T545 = R546;
  assign io_yout_4 = yout_4;
  assign yout_4 = T547;
  assign T547 = T612 + T548;
  assign T548 = R549;
  assign T550 = T1178;
  assign T1178 = T551[5'h11:1'h0];
  assign T551 = $signed(T552) >>> 4'he;
  assign T552 = $signed(T554) * $signed(T553);
  assign T553 = 18'h8000;
  assign T554 = T555;
  assign T555 = T1179;
  assign T1179 = T556[5'h11:1'h0];
  assign T556 = $signed(T557) >>> 4'he;
  assign T557 = $signed(T559) * $signed(T558);
  assign T558 = io_lbda;
  assign T559 = T560;
  assign T560 = T561;
  assign T561 = T566 - T562;
  assign T562 = R563;
  assign T566 = R567;
  assign T569 = T609 ? 18'h8000 : T570;
  assign T570 = T606 ? 18'h38000 : T571;
  assign T571 = T572;
  assign T572 = T574 + T573;
  assign T573 = R565;
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T579 - T577;
  assign T577 = R578;
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = T589 + T582;
  assign T582 = T583;
  assign T583 = T1180;
  assign T1180 = T584[5'h11:1'h0];
  assign T584 = $signed(T585) >>> 4'he;
  assign T585 = $signed(T587) * $signed(T586);
  assign T586 = R33;
  assign T587 = R588;
  assign T589 = T590;
  assign T590 = T591;
  assign T591 = T599 + T592;
  assign T592 = T593;
  assign T593 = T1181;
  assign T1181 = T594[5'h11:1'h0];
  assign T594 = $signed(T595) >>> 4'he;
  assign T595 = $signed(T597) * $signed(T596);
  assign T596 = R46;
  assign T597 = R598;
  assign T599 = T600;
  assign T600 = T1182;
  assign T1182 = T601[5'h11:1'h0];
  assign T601 = $signed(T602) >>> 4'he;
  assign T602 = $signed(T604) * $signed(T603);
  assign T603 = R56;
  assign T604 = R605;
  assign T606 = $signed(T608) < $signed(T607);
  assign T607 = 18'h38000;
  assign T608 = T571;
  assign T609 = $signed(T611) < $signed(T610);
  assign T610 = T571;
  assign T611 = 18'h8000;
  assign T612 = R613;
  assign io_yout_5 = yout_5;
  assign yout_5 = T614;
  assign T614 = T679 + T615;
  assign T615 = R616;
  assign T617 = T1183;
  assign T1183 = T618[5'h11:1'h0];
  assign T618 = $signed(T619) >>> 4'he;
  assign T619 = $signed(T621) * $signed(T620);
  assign T620 = 18'h8000;
  assign T621 = T622;
  assign T622 = T1184;
  assign T1184 = T623[5'h11:1'h0];
  assign T623 = $signed(T624) >>> 4'he;
  assign T624 = $signed(T626) * $signed(T625);
  assign T625 = io_lbda;
  assign T626 = T627;
  assign T627 = T628;
  assign T628 = T633 - T629;
  assign T629 = R630;
  assign T633 = R634;
  assign T636 = T676 ? 18'h8000 : T637;
  assign T637 = T673 ? 18'h38000 : T638;
  assign T638 = T639;
  assign T639 = T641 + T640;
  assign T640 = R632;
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = T646 - T644;
  assign T644 = R645;
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T656 + T649;
  assign T649 = T650;
  assign T650 = T1185;
  assign T1185 = T651[5'h11:1'h0];
  assign T651 = $signed(T652) >>> 4'he;
  assign T652 = $signed(T654) * $signed(T653);
  assign T653 = R33;
  assign T654 = R655;
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T666 + T659;
  assign T659 = T660;
  assign T660 = T1186;
  assign T1186 = T661[5'h11:1'h0];
  assign T661 = $signed(T662) >>> 4'he;
  assign T662 = $signed(T664) * $signed(T663);
  assign T663 = R46;
  assign T664 = R665;
  assign T666 = T667;
  assign T667 = T1187;
  assign T1187 = T668[5'h11:1'h0];
  assign T668 = $signed(T669) >>> 4'he;
  assign T669 = $signed(T671) * $signed(T670);
  assign T670 = R56;
  assign T671 = R672;
  assign T673 = $signed(T675) < $signed(T674);
  assign T674 = 18'h38000;
  assign T675 = T638;
  assign T676 = $signed(T678) < $signed(T677);
  assign T677 = T638;
  assign T678 = 18'h8000;
  assign T679 = R680;
  assign io_yout_6 = yout_6;
  assign yout_6 = T681;
  assign T681 = T746 + T682;
  assign T682 = R683;
  assign T684 = T1188;
  assign T1188 = T685[5'h11:1'h0];
  assign T685 = $signed(T686) >>> 4'he;
  assign T686 = $signed(T688) * $signed(T687);
  assign T687 = 18'h8000;
  assign T688 = T689;
  assign T689 = T1189;
  assign T1189 = T690[5'h11:1'h0];
  assign T690 = $signed(T691) >>> 4'he;
  assign T691 = $signed(T693) * $signed(T692);
  assign T692 = io_lbda;
  assign T693 = T694;
  assign T694 = T695;
  assign T695 = T700 - T696;
  assign T696 = R697;
  assign T700 = R701;
  assign T703 = T743 ? 18'h8000 : T704;
  assign T704 = T740 ? 18'h38000 : T705;
  assign T705 = T706;
  assign T706 = T708 + T707;
  assign T707 = R699;
  assign T708 = T709;
  assign T709 = T710;
  assign T710 = T713 - T711;
  assign T711 = R712;
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = T723 + T716;
  assign T716 = T717;
  assign T717 = T1190;
  assign T1190 = T718[5'h11:1'h0];
  assign T718 = $signed(T719) >>> 4'he;
  assign T719 = $signed(T721) * $signed(T720);
  assign T720 = R33;
  assign T721 = R722;
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = T733 + T726;
  assign T726 = T727;
  assign T727 = T1191;
  assign T1191 = T728[5'h11:1'h0];
  assign T728 = $signed(T729) >>> 4'he;
  assign T729 = $signed(T731) * $signed(T730);
  assign T730 = R46;
  assign T731 = R732;
  assign T733 = T734;
  assign T734 = T1192;
  assign T1192 = T735[5'h11:1'h0];
  assign T735 = $signed(T736) >>> 4'he;
  assign T736 = $signed(T738) * $signed(T737);
  assign T737 = R56;
  assign T738 = R739;
  assign T740 = $signed(T742) < $signed(T741);
  assign T741 = 18'h38000;
  assign T742 = T705;
  assign T743 = $signed(T745) < $signed(T744);
  assign T744 = T705;
  assign T745 = 18'h8000;
  assign T746 = R747;
  assign io_yout_7 = yout_7;
  assign yout_7 = T748;
  assign T748 = T813 + T749;
  assign T749 = R750;
  assign T751 = T1193;
  assign T1193 = T752[5'h11:1'h0];
  assign T752 = $signed(T753) >>> 4'he;
  assign T753 = $signed(T755) * $signed(T754);
  assign T754 = 18'h8000;
  assign T755 = T756;
  assign T756 = T1194;
  assign T1194 = T757[5'h11:1'h0];
  assign T757 = $signed(T758) >>> 4'he;
  assign T758 = $signed(T760) * $signed(T759);
  assign T759 = io_lbda;
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T767 - T763;
  assign T763 = R764;
  assign T767 = R768;
  assign T770 = T810 ? 18'h8000 : T771;
  assign T771 = T807 ? 18'h38000 : T772;
  assign T772 = T773;
  assign T773 = T775 + T774;
  assign T774 = R766;
  assign T775 = T776;
  assign T776 = T777;
  assign T777 = T780 - T778;
  assign T778 = R779;
  assign T780 = T781;
  assign T781 = T782;
  assign T782 = T790 + T783;
  assign T783 = T784;
  assign T784 = T1195;
  assign T1195 = T785[5'h11:1'h0];
  assign T785 = $signed(T786) >>> 4'he;
  assign T786 = $signed(T788) * $signed(T787);
  assign T787 = R33;
  assign T788 = R789;
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T800 + T793;
  assign T793 = T794;
  assign T794 = T1196;
  assign T1196 = T795[5'h11:1'h0];
  assign T795 = $signed(T796) >>> 4'he;
  assign T796 = $signed(T798) * $signed(T797);
  assign T797 = R46;
  assign T798 = R799;
  assign T800 = T801;
  assign T801 = T1197;
  assign T1197 = T802[5'h11:1'h0];
  assign T802 = $signed(T803) >>> 4'he;
  assign T803 = $signed(T805) * $signed(T804);
  assign T804 = R56;
  assign T805 = R806;
  assign T807 = $signed(T809) < $signed(T808);
  assign T808 = 18'h38000;
  assign T809 = T772;
  assign T810 = $signed(T812) < $signed(T811);
  assign T811 = T772;
  assign T812 = 18'h8000;
  assign T813 = R814;
  assign io_yout_8 = yout_8;
  assign yout_8 = T815;
  assign T815 = T880 + T816;
  assign T816 = R817;
  assign T818 = T1198;
  assign T1198 = T819[5'h11:1'h0];
  assign T819 = $signed(T820) >>> 4'he;
  assign T820 = $signed(T822) * $signed(T821);
  assign T821 = 18'h8000;
  assign T822 = T823;
  assign T823 = T1199;
  assign T1199 = T824[5'h11:1'h0];
  assign T824 = $signed(T825) >>> 4'he;
  assign T825 = $signed(T827) * $signed(T826);
  assign T826 = io_lbda;
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = T834 - T830;
  assign T830 = R831;
  assign T834 = R835;
  assign T837 = T877 ? 18'h8000 : T838;
  assign T838 = T874 ? 18'h38000 : T839;
  assign T839 = T840;
  assign T840 = T842 + T841;
  assign T841 = R833;
  assign T842 = T843;
  assign T843 = T844;
  assign T844 = T847 - T845;
  assign T845 = R846;
  assign T847 = T848;
  assign T848 = T849;
  assign T849 = T857 + T850;
  assign T850 = T851;
  assign T851 = T1200;
  assign T1200 = T852[5'h11:1'h0];
  assign T852 = $signed(T853) >>> 4'he;
  assign T853 = $signed(T855) * $signed(T854);
  assign T854 = R33;
  assign T855 = R856;
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = T867 + T860;
  assign T860 = T861;
  assign T861 = T1201;
  assign T1201 = T862[5'h11:1'h0];
  assign T862 = $signed(T863) >>> 4'he;
  assign T863 = $signed(T865) * $signed(T864);
  assign T864 = R46;
  assign T865 = R866;
  assign T867 = T868;
  assign T868 = T1202;
  assign T1202 = T869[5'h11:1'h0];
  assign T869 = $signed(T870) >>> 4'he;
  assign T870 = $signed(T872) * $signed(T871);
  assign T871 = R56;
  assign T872 = R873;
  assign T874 = $signed(T876) < $signed(T875);
  assign T875 = 18'h38000;
  assign T876 = T839;
  assign T877 = $signed(T879) < $signed(T878);
  assign T878 = T839;
  assign T879 = 18'h8000;
  assign T880 = R881;
  assign io_yout_9 = yout_9;
  assign yout_9 = T882;
  assign T882 = T947 + T883;
  assign T883 = R884;
  assign T885 = T1203;
  assign T1203 = T886[5'h11:1'h0];
  assign T886 = $signed(T887) >>> 4'he;
  assign T887 = $signed(T889) * $signed(T888);
  assign T888 = 18'h8000;
  assign T889 = T890;
  assign T890 = T1204;
  assign T1204 = T891[5'h11:1'h0];
  assign T891 = $signed(T892) >>> 4'he;
  assign T892 = $signed(T894) * $signed(T893);
  assign T893 = io_lbda;
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T901 - T897;
  assign T897 = R898;
  assign T901 = R902;
  assign T904 = T944 ? 18'h8000 : T905;
  assign T905 = T941 ? 18'h38000 : T906;
  assign T906 = T907;
  assign T907 = T909 + T908;
  assign T908 = R900;
  assign T909 = T910;
  assign T910 = T911;
  assign T911 = T914 - T912;
  assign T912 = R913;
  assign T914 = T915;
  assign T915 = T916;
  assign T916 = T924 + T917;
  assign T917 = T918;
  assign T918 = T1205;
  assign T1205 = T919[5'h11:1'h0];
  assign T919 = $signed(T920) >>> 4'he;
  assign T920 = $signed(T922) * $signed(T921);
  assign T921 = R33;
  assign T922 = R923;
  assign T924 = T925;
  assign T925 = T926;
  assign T926 = T934 + T927;
  assign T927 = T928;
  assign T928 = T1206;
  assign T1206 = T929[5'h11:1'h0];
  assign T929 = $signed(T930) >>> 4'he;
  assign T930 = $signed(T932) * $signed(T931);
  assign T931 = R46;
  assign T932 = R933;
  assign T934 = T935;
  assign T935 = T1207;
  assign T1207 = T936[5'h11:1'h0];
  assign T936 = $signed(T937) >>> 4'he;
  assign T937 = $signed(T939) * $signed(T938);
  assign T938 = R56;
  assign T939 = R940;
  assign T941 = $signed(T943) < $signed(T942);
  assign T942 = 18'h38000;
  assign T943 = T906;
  assign T944 = $signed(T946) < $signed(T945);
  assign T945 = T906;
  assign T946 = 18'h8000;
  assign T947 = R948;
  assign io_yout_10 = yout_10;
  assign yout_10 = T949;
  assign T949 = T1014 + T950;
  assign T950 = R951;
  assign T952 = T1208;
  assign T1208 = T953[5'h11:1'h0];
  assign T953 = $signed(T954) >>> 4'he;
  assign T954 = $signed(T956) * $signed(T955);
  assign T955 = 18'h8000;
  assign T956 = T957;
  assign T957 = T1209;
  assign T1209 = T958[5'h11:1'h0];
  assign T958 = $signed(T959) >>> 4'he;
  assign T959 = $signed(T961) * $signed(T960);
  assign T960 = io_lbda;
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = T968 - T964;
  assign T964 = R965;
  assign T968 = R969;
  assign T971 = T1011 ? 18'h8000 : T972;
  assign T972 = T1008 ? 18'h38000 : T973;
  assign T973 = T974;
  assign T974 = T976 + T975;
  assign T975 = R967;
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T981 - T979;
  assign T979 = R980;
  assign T981 = T982;
  assign T982 = T983;
  assign T983 = T991 + T984;
  assign T984 = T985;
  assign T985 = T1210;
  assign T1210 = T986[5'h11:1'h0];
  assign T986 = $signed(T987) >>> 4'he;
  assign T987 = $signed(T989) * $signed(T988);
  assign T988 = R33;
  assign T989 = R990;
  assign T991 = T992;
  assign T992 = T993;
  assign T993 = T1001 + T994;
  assign T994 = T995;
  assign T995 = T1211;
  assign T1211 = T996[5'h11:1'h0];
  assign T996 = $signed(T997) >>> 4'he;
  assign T997 = $signed(T999) * $signed(T998);
  assign T998 = R46;
  assign T999 = R1000;
  assign T1001 = T1002;
  assign T1002 = T1212;
  assign T1212 = T1003[5'h11:1'h0];
  assign T1003 = $signed(T1004) >>> 4'he;
  assign T1004 = $signed(T1006) * $signed(T1005);
  assign T1005 = R56;
  assign T1006 = R1007;
  assign T1008 = $signed(T1010) < $signed(T1009);
  assign T1009 = 18'h38000;
  assign T1010 = T973;
  assign T1011 = $signed(T1013) < $signed(T1012);
  assign T1012 = T973;
  assign T1013 = 18'h8000;
  assign T1014 = R1015;
  assign io_yout_11 = yout_11;
  assign yout_11 = T1016;
  assign T1016 = T1081 + T1017;
  assign T1017 = R1018;
  assign T1019 = T1213;
  assign T1213 = T1020[5'h11:1'h0];
  assign T1020 = $signed(T1021) >>> 4'he;
  assign T1021 = $signed(T1023) * $signed(T1022);
  assign T1022 = 18'h8000;
  assign T1023 = T1024;
  assign T1024 = T1214;
  assign T1214 = T1025[5'h11:1'h0];
  assign T1025 = $signed(T1026) >>> 4'he;
  assign T1026 = $signed(T1028) * $signed(T1027);
  assign T1027 = io_lbda;
  assign T1028 = T1029;
  assign T1029 = T1030;
  assign T1030 = T1035 - T1031;
  assign T1031 = R1032;
  assign T1035 = R1036;
  assign T1038 = T1078 ? 18'h8000 : T1039;
  assign T1039 = T1075 ? 18'h38000 : T1040;
  assign T1040 = T1041;
  assign T1041 = T1043 + T1042;
  assign T1042 = R1034;
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = T1048 - T1046;
  assign T1046 = R1047;
  assign T1048 = T1049;
  assign T1049 = T1050;
  assign T1050 = T1058 + T1051;
  assign T1051 = T1052;
  assign T1052 = T1215;
  assign T1215 = T1053[5'h11:1'h0];
  assign T1053 = $signed(T1054) >>> 4'he;
  assign T1054 = $signed(T1056) * $signed(T1055);
  assign T1055 = R33;
  assign T1056 = R1057;
  assign T1058 = T1059;
  assign T1059 = T1060;
  assign T1060 = T1068 + T1061;
  assign T1061 = T1062;
  assign T1062 = T1216;
  assign T1216 = T1063[5'h11:1'h0];
  assign T1063 = $signed(T1064) >>> 4'he;
  assign T1064 = $signed(T1066) * $signed(T1065);
  assign T1065 = R46;
  assign T1066 = R1067;
  assign T1068 = T1069;
  assign T1069 = T1217;
  assign T1217 = T1070[5'h11:1'h0];
  assign T1070 = $signed(T1071) >>> 4'he;
  assign T1071 = $signed(T1073) * $signed(T1072);
  assign T1072 = R56;
  assign T1073 = R1074;
  assign T1075 = $signed(T1077) < $signed(T1076);
  assign T1076 = 18'h38000;
  assign T1077 = T1040;
  assign T1078 = $signed(T1080) < $signed(T1079);
  assign T1079 = T1040;
  assign T1080 = 18'h8000;
  assign T1081 = R1082;
  assign io_xout_0 = xout_0;
  assign xout_0 = T1083;
  assign T1083 = T1098 + T1084;
  assign T1084 = R1085;
  assign T1086 = T1218;
  assign T1218 = T1087[5'h11:1'h0];
  assign T1087 = $signed(T1088) >>> 4'he;
  assign T1088 = $signed(T1090) * $signed(T1089);
  assign T1089 = io_lbda;
  assign T1090 = T1091;
  assign T1091 = T1092;
  assign T1092 = T1097 - T1093;
  assign T1093 = R1094;
  assign T1097 = R93;
  assign T1098 = R1099;
  assign io_xout_1 = xout_1;
  assign xout_1 = T1100;
  assign T1100 = T1115 + T1101;
  assign T1101 = R1102;
  assign T1103 = T1219;
  assign T1219 = T1104[5'h11:1'h0];
  assign T1104 = $signed(T1105) >>> 4'he;
  assign T1105 = $signed(T1107) * $signed(T1106);
  assign T1106 = io_lbda;
  assign T1107 = T1108;
  assign T1108 = T1109;
  assign T1109 = T1114 - T1110;
  assign T1110 = R1111;
  assign T1114 = R85;
  assign T1115 = R1116;
  assign io_xout_2 = xout_2;
  assign xout_2 = T1117;
  assign T1117 = T1132 + T1118;
  assign T1118 = R1119;
  assign T1120 = T1220;
  assign T1220 = T1121[5'h11:1'h0];
  assign T1121 = $signed(T1122) >>> 4'he;
  assign T1122 = $signed(T1124) * $signed(T1123);
  assign T1123 = io_lbda;
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1131 - T1127;
  assign T1127 = R1128;
  assign T1131 = R74;
  assign T1132 = R1133;
  XNetModule XNetModule(
       .io_x_2( io_x_2 ),
       .io_x_1( io_x_1 ),
       .io_x_0( io_x_0 ),
       .io_y_11( io_y_11 ),
       .io_y_10( io_y_10 ),
       .io_y_9( io_y_9 ),
       .io_y_8( io_y_8 ),
       .io_y_7( io_y_7 ),
       .io_y_6( io_y_6 ),
       .io_y_5( io_y_5 ),
       .io_y_4( io_y_4 ),
       .io_y_3( io_y_3 ),
       .io_y_2( io_y_2 ),
       .io_y_1( io_y_1 ),
       .io_y_0( io_y_0 ),
       .io_z_2( io_z_2 ),
       .io_z_1( io_z_1 ),
       .io_z_0( io_z_0 ),
       .io_a_11_2( io_a_11_2 ),
       .io_a_11_1( io_a_11_1 ),
       .io_a_11_0( io_a_11_0 ),
       .io_a_10_2( io_a_10_2 ),
       .io_a_10_1( io_a_10_1 ),
       .io_a_10_0( io_a_10_0 ),
       .io_a_9_2( io_a_9_2 ),
       .io_a_9_1( io_a_9_1 ),
       .io_a_9_0( io_a_9_0 ),
       .io_a_8_2( io_a_8_2 ),
       .io_a_8_1( io_a_8_1 ),
       .io_a_8_0( io_a_8_0 ),
       .io_a_7_2( io_a_7_2 ),
       .io_a_7_1( io_a_7_1 ),
       .io_a_7_0( io_a_7_0 ),
       .io_a_6_2( io_a_6_2 ),
       .io_a_6_1( io_a_6_1 ),
       .io_a_6_0( io_a_6_0 ),
       .io_a_5_2( io_a_5_2 ),
       .io_a_5_1( io_a_5_1 ),
       .io_a_5_0( io_a_5_0 ),
       .io_a_4_2( io_a_4_2 ),
       .io_a_4_1( io_a_4_1 ),
       .io_a_4_0( io_a_4_0 ),
       .io_a_3_2( io_a_3_2 ),
       .io_a_3_1( io_a_3_1 ),
       .io_a_3_0( io_a_3_0 ),
       .io_a_2_2( io_a_2_2 ),
       .io_a_2_1( io_a_2_1 ),
       .io_a_2_0( io_a_2_0 ),
       .io_a_1_2( io_a_1_2 ),
       .io_a_1_1( io_a_1_1 ),
       .io_a_1_0( io_a_1_0 ),
       .io_a_0_2( io_a_0_2 ),
       .io_a_0_1( io_a_0_1 ),
       .io_a_0_0( io_a_0_0 ),
       .io_c_2_2( io_c_2_2 ),
       .io_c_2_1( io_c_2_1 ),
       .io_c_2_0( io_c_2_0 ),
       .io_c_1_2( io_c_1_2 ),
       .io_c_1_1( io_c_1_1 ),
       .io_c_1_0( io_c_1_0 ),
       .io_c_0_2( io_c_0_2 ),
       .io_c_0_1( io_c_0_1 ),
       .io_c_0_0( io_c_0_0 ),
       .io_o_2( XNetModule_io_o_2 ),
       .io_o_1( XNetModule_io_o_1 ),
       .io_o_0( XNetModule_io_o_0 )
  );

  always @(posedge clk) begin
    R2 <= T3;
    if(T63) begin
      R16 <= 18'h8000;
    end else if(T60) begin
      R16 <= 18'h38000;
    end else begin
      R16 <= T19;
    end
    R22 <= R23;
    R23 <= io_z_0;
    R32 <= R33;
    R33 <= XNetModule_io_o_2;
    R35 <= R36;
    R36 <= io_c_0_2;
    R45 <= R46;
    R46 <= XNetModule_io_o_1;
    R48 <= R49;
    R49 <= io_c_0_1;
    R55 <= R56;
    R56 <= XNetModule_io_o_0;
    R58 <= R59;
    R59 <= io_c_0_0;
    R74 <= R32;
    R76 <= R35;
    R85 <= R45;
    R87 <= R48;
    R93 <= R55;
    R95 <= R58;
    R97 <= R98;
    R98 <= R22;
    R101 <= T102;
    if(T156) begin
      R115 <= 18'h8000;
    end else if(T153) begin
      R115 <= 18'h38000;
    end else begin
      R115 <= T118;
    end
    R121 <= R122;
    R122 <= io_z_1;
    R132 <= R133;
    R133 <= io_c_1_2;
    R143 <= R144;
    R144 <= io_c_1_1;
    R151 <= R152;
    R152 <= io_c_1_0;
    R168 <= R132;
    R178 <= R143;
    R185 <= R151;
    R187 <= R188;
    R188 <= R121;
    R191 <= T192;
    if(T246) begin
      R205 <= 18'h8000;
    end else if(T243) begin
      R205 <= 18'h38000;
    end else begin
      R205 <= T208;
    end
    R211 <= R212;
    R212 <= io_z_2;
    R222 <= R223;
    R223 <= io_c_2_2;
    R233 <= R234;
    R234 <= io_c_2_1;
    R241 <= R242;
    R242 <= io_c_2_0;
    R258 <= R222;
    R268 <= R233;
    R275 <= R241;
    R277 <= R278;
    R278 <= R211;
    R281 <= T282;
    R295 <= R296;
    R296 <= R297;
    R297 <= io_y_0;
    R299 <= R300;
    if(T341) begin
      R300 <= 18'h8000;
    end else if(T338) begin
      R300 <= 18'h38000;
    end else begin
      R300 <= T303;
    end
    R310 <= io_b_0;
    R320 <= io_a_0_2;
    R330 <= io_a_0_1;
    R337 <= io_a_0_0;
    R345 <= R295;
    R348 <= T349;
    R362 <= R363;
    R363 <= R364;
    R364 <= io_y_1;
    R366 <= R367;
    if(T408) begin
      R367 <= 18'h8000;
    end else if(T405) begin
      R367 <= 18'h38000;
    end else begin
      R367 <= T370;
    end
    R377 <= io_b_1;
    R387 <= io_a_1_2;
    R397 <= io_a_1_1;
    R404 <= io_a_1_0;
    R412 <= R362;
    R415 <= T416;
    R429 <= R430;
    R430 <= R431;
    R431 <= io_y_2;
    R433 <= R434;
    if(T475) begin
      R434 <= 18'h8000;
    end else if(T472) begin
      R434 <= 18'h38000;
    end else begin
      R434 <= T437;
    end
    R444 <= io_b_2;
    R454 <= io_a_2_2;
    R464 <= io_a_2_1;
    R471 <= io_a_2_0;
    R479 <= R429;
    R482 <= T483;
    R496 <= R497;
    R497 <= R498;
    R498 <= io_y_3;
    R500 <= R501;
    if(T542) begin
      R501 <= 18'h8000;
    end else if(T539) begin
      R501 <= 18'h38000;
    end else begin
      R501 <= T504;
    end
    R511 <= io_b_3;
    R521 <= io_a_3_2;
    R531 <= io_a_3_1;
    R538 <= io_a_3_0;
    R546 <= R496;
    R549 <= T550;
    R563 <= R564;
    R564 <= R565;
    R565 <= io_y_4;
    R567 <= R568;
    if(T609) begin
      R568 <= 18'h8000;
    end else if(T606) begin
      R568 <= 18'h38000;
    end else begin
      R568 <= T571;
    end
    R578 <= io_b_4;
    R588 <= io_a_4_2;
    R598 <= io_a_4_1;
    R605 <= io_a_4_0;
    R613 <= R563;
    R616 <= T617;
    R630 <= R631;
    R631 <= R632;
    R632 <= io_y_5;
    R634 <= R635;
    if(T676) begin
      R635 <= 18'h8000;
    end else if(T673) begin
      R635 <= 18'h38000;
    end else begin
      R635 <= T638;
    end
    R645 <= io_b_5;
    R655 <= io_a_5_2;
    R665 <= io_a_5_1;
    R672 <= io_a_5_0;
    R680 <= R630;
    R683 <= T684;
    R697 <= R698;
    R698 <= R699;
    R699 <= io_y_6;
    R701 <= R702;
    if(T743) begin
      R702 <= 18'h8000;
    end else if(T740) begin
      R702 <= 18'h38000;
    end else begin
      R702 <= T705;
    end
    R712 <= io_b_6;
    R722 <= io_a_6_2;
    R732 <= io_a_6_1;
    R739 <= io_a_6_0;
    R747 <= R697;
    R750 <= T751;
    R764 <= R765;
    R765 <= R766;
    R766 <= io_y_7;
    R768 <= R769;
    if(T810) begin
      R769 <= 18'h8000;
    end else if(T807) begin
      R769 <= 18'h38000;
    end else begin
      R769 <= T772;
    end
    R779 <= io_b_7;
    R789 <= io_a_7_2;
    R799 <= io_a_7_1;
    R806 <= io_a_7_0;
    R814 <= R764;
    R817 <= T818;
    R831 <= R832;
    R832 <= R833;
    R833 <= io_y_8;
    R835 <= R836;
    if(T877) begin
      R836 <= 18'h8000;
    end else if(T874) begin
      R836 <= 18'h38000;
    end else begin
      R836 <= T839;
    end
    R846 <= io_b_8;
    R856 <= io_a_8_2;
    R866 <= io_a_8_1;
    R873 <= io_a_8_0;
    R881 <= R831;
    R884 <= T885;
    R898 <= R899;
    R899 <= R900;
    R900 <= io_y_9;
    R902 <= R903;
    if(T944) begin
      R903 <= 18'h8000;
    end else if(T941) begin
      R903 <= 18'h38000;
    end else begin
      R903 <= T906;
    end
    R913 <= io_b_9;
    R923 <= io_a_9_2;
    R933 <= io_a_9_1;
    R940 <= io_a_9_0;
    R948 <= R898;
    R951 <= T952;
    R965 <= R966;
    R966 <= R967;
    R967 <= io_y_10;
    R969 <= R970;
    if(T1011) begin
      R970 <= 18'h8000;
    end else if(T1008) begin
      R970 <= 18'h38000;
    end else begin
      R970 <= T973;
    end
    R980 <= io_b_10;
    R990 <= io_a_10_2;
    R1000 <= io_a_10_1;
    R1007 <= io_a_10_0;
    R1015 <= R965;
    R1018 <= T1019;
    R1032 <= R1033;
    R1033 <= R1034;
    R1034 <= io_y_11;
    R1036 <= R1037;
    if(T1078) begin
      R1037 <= 18'h8000;
    end else if(T1075) begin
      R1037 <= 18'h38000;
    end else begin
      R1037 <= T1040;
    end
    R1047 <= io_b_11;
    R1057 <= io_a_11_2;
    R1067 <= io_a_11_1;
    R1074 <= io_a_11_0;
    R1082 <= R1032;
    R1085 <= T1086;
    R1094 <= R1095;
    R1095 <= R1096;
    R1096 <= io_x_0;
    R1099 <= R1094;
    R1102 <= T1103;
    R1111 <= R1112;
    R1112 <= R1113;
    R1113 <= io_x_1;
    R1116 <= R1111;
    R1119 <= T1120;
    R1128 <= R1129;
    R1129 <= R1130;
    R1130 <= io_x_2;
    R1133 <= R1128;
  end
endmodule

module NN1ShiftTop(input clk, input reset,
    input [17:0] io_x,
    input [17:0] io_y,
    input [17:0] io_z,
    input [17:0] io_b,
    input [17:0] io_a,
    input [17:0] io_c,
    input [17:0] io_lbda,
    output[17:0] io_xout,
    output[17:0] io_yout,
    output[17:0] io_zout
);

  reg [17:0] cShift_0_0;
  wire[17:0] T60;
  reg [17:0] cShift_1_0;
  wire[17:0] T61;
  reg [17:0] cShift_2_0;
  wire[17:0] T62;
  reg [17:0] cShift_0_1;
  wire[17:0] T63;
  reg [17:0] cShift_1_1;
  wire[17:0] T64;
  reg [17:0] cShift_2_1;
  wire[17:0] T65;
  reg [17:0] cShift_0_2;
  wire[17:0] T66;
  reg [17:0] cShift_1_2;
  wire[17:0] T67;
  reg [17:0] cShift_2_2;
  wire[17:0] T68;
  reg [17:0] aShift_0_0;
  wire[17:0] T69;
  reg [17:0] aShift_1_0;
  wire[17:0] T70;
  reg [17:0] aShift_2_0;
  wire[17:0] T71;
  reg [17:0] aShift_3_0;
  wire[17:0] T72;
  reg [17:0] aShift_4_0;
  wire[17:0] T73;
  reg [17:0] aShift_5_0;
  wire[17:0] T74;
  reg [17:0] aShift_6_0;
  wire[17:0] T75;
  reg [17:0] aShift_7_0;
  wire[17:0] T76;
  reg [17:0] aShift_8_0;
  wire[17:0] T77;
  reg [17:0] aShift_9_0;
  wire[17:0] T78;
  reg [17:0] aShift_10_0;
  wire[17:0] T79;
  reg [17:0] aShift_11_0;
  wire[17:0] T80;
  reg [17:0] aShift_0_1;
  wire[17:0] T81;
  reg [17:0] aShift_1_1;
  wire[17:0] T82;
  reg [17:0] aShift_2_1;
  wire[17:0] T83;
  reg [17:0] aShift_3_1;
  wire[17:0] T84;
  reg [17:0] aShift_4_1;
  wire[17:0] T85;
  reg [17:0] aShift_5_1;
  wire[17:0] T86;
  reg [17:0] aShift_6_1;
  wire[17:0] T87;
  reg [17:0] aShift_7_1;
  wire[17:0] T88;
  reg [17:0] aShift_8_1;
  wire[17:0] T89;
  reg [17:0] aShift_9_1;
  wire[17:0] T90;
  reg [17:0] aShift_10_1;
  wire[17:0] T91;
  reg [17:0] aShift_11_1;
  wire[17:0] T92;
  reg [17:0] aShift_0_2;
  wire[17:0] T93;
  reg [17:0] aShift_1_2;
  wire[17:0] T94;
  reg [17:0] aShift_2_2;
  wire[17:0] T95;
  reg [17:0] aShift_3_2;
  wire[17:0] T96;
  reg [17:0] aShift_4_2;
  wire[17:0] T97;
  reg [17:0] aShift_5_2;
  wire[17:0] T98;
  reg [17:0] aShift_6_2;
  wire[17:0] T99;
  reg [17:0] aShift_7_2;
  wire[17:0] T100;
  reg [17:0] aShift_8_2;
  wire[17:0] T101;
  reg [17:0] aShift_9_2;
  wire[17:0] T102;
  reg [17:0] aShift_10_2;
  wire[17:0] T103;
  reg [17:0] aShift_11_2;
  wire[17:0] T104;
  reg [17:0] bShift_0;
  wire[17:0] T105;
  reg [17:0] bShift_1;
  wire[17:0] T106;
  reg [17:0] bShift_2;
  wire[17:0] T107;
  reg [17:0] bShift_3;
  wire[17:0] T108;
  reg [17:0] bShift_4;
  wire[17:0] T109;
  reg [17:0] bShift_5;
  wire[17:0] T110;
  reg [17:0] bShift_6;
  wire[17:0] T111;
  reg [17:0] bShift_7;
  wire[17:0] T112;
  reg [17:0] bShift_8;
  wire[17:0] T113;
  reg [17:0] bShift_9;
  wire[17:0] T114;
  reg [17:0] bShift_10;
  wire[17:0] T115;
  reg [17:0] bShift_11;
  wire[17:0] T116;
  reg [17:0] zShift_0;
  wire[17:0] T117;
  reg [17:0] zShift_1;
  wire[17:0] T118;
  reg [17:0] zShift_2;
  wire[17:0] T119;
  reg [17:0] yShift_0;
  wire[17:0] T120;
  reg [17:0] yShift_1;
  wire[17:0] T121;
  reg [17:0] yShift_2;
  wire[17:0] T122;
  reg [17:0] yShift_3;
  wire[17:0] T123;
  reg [17:0] yShift_4;
  wire[17:0] T124;
  reg [17:0] yShift_5;
  wire[17:0] T125;
  reg [17:0] yShift_6;
  wire[17:0] T126;
  reg [17:0] yShift_7;
  wire[17:0] T127;
  reg [17:0] yShift_8;
  wire[17:0] T128;
  reg [17:0] yShift_9;
  wire[17:0] T129;
  reg [17:0] yShift_10;
  wire[17:0] T130;
  reg [17:0] yShift_11;
  wire[17:0] T131;
  reg [17:0] xShift_0;
  wire[17:0] T132;
  reg [17:0] xShift_1;
  wire[17:0] T133;
  reg [17:0] xShift_2;
  wire[17:0] T134;
  reg [17:0] nnzout;
  wire[17:0] T0;
  wire[17:0] T1;
  wire[17:0] T2;
  wire[17:0] T3;
  wire[17:0] T4;
  wire[17:0] T5;
  wire[17:0] T6;
  wire[17:0] T7;
  reg [17:0] nnyout;
  wire[17:0] T8;
  wire[17:0] T9;
  wire[17:0] T10;
  wire[17:0] T11;
  wire[17:0] T12;
  wire[17:0] T13;
  wire[17:0] T14;
  wire[17:0] T15;
  wire[17:0] T16;
  wire[17:0] T17;
  wire[17:0] T18;
  wire[17:0] T19;
  wire[17:0] T20;
  wire[17:0] T21;
  wire[17:0] T22;
  wire[17:0] T23;
  wire[17:0] T24;
  wire[17:0] T25;
  wire[17:0] T26;
  wire[17:0] T27;
  wire[17:0] T28;
  wire[17:0] T29;
  wire[17:0] T30;
  wire[17:0] T31;
  wire[17:0] T32;
  wire[17:0] T33;
  wire[17:0] T34;
  wire[17:0] T35;
  wire[17:0] T36;
  wire[17:0] T37;
  wire[17:0] T38;
  wire[17:0] T39;
  wire[17:0] T40;
  wire[17:0] T41;
  wire[17:0] T42;
  wire[17:0] T43;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[17:0] T46;
  wire[17:0] T47;
  wire[17:0] T48;
  wire[17:0] T49;
  wire[17:0] T50;
  wire[17:0] T51;
  reg [17:0] nnxout;
  wire[17:0] T52;
  wire[17:0] T53;
  wire[17:0] T54;
  wire[17:0] T55;
  wire[17:0] T56;
  wire[17:0] T57;
  wire[17:0] T58;
  wire[17:0] T59;
  wire[17:0] nnTop_io_xout_2;
  wire[17:0] nnTop_io_xout_1;
  wire[17:0] nnTop_io_xout_0;
  wire[17:0] nnTop_io_yout_11;
  wire[17:0] nnTop_io_yout_10;
  wire[17:0] nnTop_io_yout_9;
  wire[17:0] nnTop_io_yout_8;
  wire[17:0] nnTop_io_yout_7;
  wire[17:0] nnTop_io_yout_6;
  wire[17:0] nnTop_io_yout_5;
  wire[17:0] nnTop_io_yout_4;
  wire[17:0] nnTop_io_yout_3;
  wire[17:0] nnTop_io_yout_2;
  wire[17:0] nnTop_io_yout_1;
  wire[17:0] nnTop_io_yout_0;
  wire[17:0] nnTop_io_zout_2;
  wire[17:0] nnTop_io_zout_1;
  wire[17:0] nnTop_io_zout_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    cShift_0_0 = {1{$random}};
    cShift_1_0 = {1{$random}};
    cShift_2_0 = {1{$random}};
    cShift_0_1 = {1{$random}};
    cShift_1_1 = {1{$random}};
    cShift_2_1 = {1{$random}};
    cShift_0_2 = {1{$random}};
    cShift_1_2 = {1{$random}};
    cShift_2_2 = {1{$random}};
    aShift_0_0 = {1{$random}};
    aShift_1_0 = {1{$random}};
    aShift_2_0 = {1{$random}};
    aShift_3_0 = {1{$random}};
    aShift_4_0 = {1{$random}};
    aShift_5_0 = {1{$random}};
    aShift_6_0 = {1{$random}};
    aShift_7_0 = {1{$random}};
    aShift_8_0 = {1{$random}};
    aShift_9_0 = {1{$random}};
    aShift_10_0 = {1{$random}};
    aShift_11_0 = {1{$random}};
    aShift_0_1 = {1{$random}};
    aShift_1_1 = {1{$random}};
    aShift_2_1 = {1{$random}};
    aShift_3_1 = {1{$random}};
    aShift_4_1 = {1{$random}};
    aShift_5_1 = {1{$random}};
    aShift_6_1 = {1{$random}};
    aShift_7_1 = {1{$random}};
    aShift_8_1 = {1{$random}};
    aShift_9_1 = {1{$random}};
    aShift_10_1 = {1{$random}};
    aShift_11_1 = {1{$random}};
    aShift_0_2 = {1{$random}};
    aShift_1_2 = {1{$random}};
    aShift_2_2 = {1{$random}};
    aShift_3_2 = {1{$random}};
    aShift_4_2 = {1{$random}};
    aShift_5_2 = {1{$random}};
    aShift_6_2 = {1{$random}};
    aShift_7_2 = {1{$random}};
    aShift_8_2 = {1{$random}};
    aShift_9_2 = {1{$random}};
    aShift_10_2 = {1{$random}};
    aShift_11_2 = {1{$random}};
    bShift_0 = {1{$random}};
    bShift_1 = {1{$random}};
    bShift_2 = {1{$random}};
    bShift_3 = {1{$random}};
    bShift_4 = {1{$random}};
    bShift_5 = {1{$random}};
    bShift_6 = {1{$random}};
    bShift_7 = {1{$random}};
    bShift_8 = {1{$random}};
    bShift_9 = {1{$random}};
    bShift_10 = {1{$random}};
    bShift_11 = {1{$random}};
    zShift_0 = {1{$random}};
    zShift_1 = {1{$random}};
    zShift_2 = {1{$random}};
    yShift_0 = {1{$random}};
    yShift_1 = {1{$random}};
    yShift_2 = {1{$random}};
    yShift_3 = {1{$random}};
    yShift_4 = {1{$random}};
    yShift_5 = {1{$random}};
    yShift_6 = {1{$random}};
    yShift_7 = {1{$random}};
    yShift_8 = {1{$random}};
    yShift_9 = {1{$random}};
    yShift_10 = {1{$random}};
    yShift_11 = {1{$random}};
    xShift_0 = {1{$random}};
    xShift_1 = {1{$random}};
    xShift_2 = {1{$random}};
    nnzout = {1{$random}};
    nnyout = {1{$random}};
    nnxout = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T60 = reset ? 18'h0 : cShift_1_0;
  assign T61 = reset ? 18'h0 : cShift_2_0;
  assign T62 = reset ? 18'h0 : io_c;
  assign T63 = reset ? 18'h0 : cShift_1_1;
  assign T64 = reset ? 18'h0 : cShift_2_1;
  assign T65 = reset ? 18'h0 : io_c;
  assign T66 = reset ? 18'h0 : cShift_1_2;
  assign T67 = reset ? 18'h0 : cShift_2_2;
  assign T68 = reset ? 18'h0 : io_c;
  assign T69 = reset ? 18'h0 : aShift_1_0;
  assign T70 = reset ? 18'h0 : aShift_2_0;
  assign T71 = reset ? 18'h0 : aShift_3_0;
  assign T72 = reset ? 18'h0 : aShift_4_0;
  assign T73 = reset ? 18'h0 : aShift_5_0;
  assign T74 = reset ? 18'h0 : aShift_6_0;
  assign T75 = reset ? 18'h0 : aShift_7_0;
  assign T76 = reset ? 18'h0 : aShift_8_0;
  assign T77 = reset ? 18'h0 : aShift_9_0;
  assign T78 = reset ? 18'h0 : aShift_10_0;
  assign T79 = reset ? 18'h0 : aShift_11_0;
  assign T80 = reset ? 18'h0 : io_a;
  assign T81 = reset ? 18'h0 : aShift_1_1;
  assign T82 = reset ? 18'h0 : aShift_2_1;
  assign T83 = reset ? 18'h0 : aShift_3_1;
  assign T84 = reset ? 18'h0 : aShift_4_1;
  assign T85 = reset ? 18'h0 : aShift_5_1;
  assign T86 = reset ? 18'h0 : aShift_6_1;
  assign T87 = reset ? 18'h0 : aShift_7_1;
  assign T88 = reset ? 18'h0 : aShift_8_1;
  assign T89 = reset ? 18'h0 : aShift_9_1;
  assign T90 = reset ? 18'h0 : aShift_10_1;
  assign T91 = reset ? 18'h0 : aShift_11_1;
  assign T92 = reset ? 18'h0 : io_a;
  assign T93 = reset ? 18'h0 : aShift_1_2;
  assign T94 = reset ? 18'h0 : aShift_2_2;
  assign T95 = reset ? 18'h0 : aShift_3_2;
  assign T96 = reset ? 18'h0 : aShift_4_2;
  assign T97 = reset ? 18'h0 : aShift_5_2;
  assign T98 = reset ? 18'h0 : aShift_6_2;
  assign T99 = reset ? 18'h0 : aShift_7_2;
  assign T100 = reset ? 18'h0 : aShift_8_2;
  assign T101 = reset ? 18'h0 : aShift_9_2;
  assign T102 = reset ? 18'h0 : aShift_10_2;
  assign T103 = reset ? 18'h0 : aShift_11_2;
  assign T104 = reset ? 18'h0 : io_a;
  assign T105 = reset ? 18'h0 : bShift_1;
  assign T106 = reset ? 18'h0 : bShift_2;
  assign T107 = reset ? 18'h0 : bShift_3;
  assign T108 = reset ? 18'h0 : bShift_4;
  assign T109 = reset ? 18'h0 : bShift_5;
  assign T110 = reset ? 18'h0 : bShift_6;
  assign T111 = reset ? 18'h0 : bShift_7;
  assign T112 = reset ? 18'h0 : bShift_8;
  assign T113 = reset ? 18'h0 : bShift_9;
  assign T114 = reset ? 18'h0 : bShift_10;
  assign T115 = reset ? 18'h0 : bShift_11;
  assign T116 = reset ? 18'h0 : io_b;
  assign T117 = reset ? 18'h0 : zShift_1;
  assign T118 = reset ? 18'h0 : zShift_2;
  assign T119 = reset ? 18'h0 : io_z;
  assign T120 = reset ? 18'h0 : yShift_1;
  assign T121 = reset ? 18'h0 : yShift_2;
  assign T122 = reset ? 18'h0 : yShift_3;
  assign T123 = reset ? 18'h0 : yShift_4;
  assign T124 = reset ? 18'h0 : yShift_5;
  assign T125 = reset ? 18'h0 : yShift_6;
  assign T126 = reset ? 18'h0 : yShift_7;
  assign T127 = reset ? 18'h0 : yShift_8;
  assign T128 = reset ? 18'h0 : yShift_9;
  assign T129 = reset ? 18'h0 : yShift_10;
  assign T130 = reset ? 18'h0 : yShift_11;
  assign T131 = reset ? 18'h0 : io_y;
  assign T132 = reset ? 18'h0 : xShift_1;
  assign T133 = reset ? 18'h0 : xShift_2;
  assign T134 = reset ? 18'h0 : io_x;
  assign io_zout = nnzout;
  assign T0 = T1;
  assign T1 = T3 + T2;
  assign T2 = nnTop_io_zout_2;
  assign T3 = T4;
  assign T4 = T5;
  assign T5 = T7 + T6;
  assign T6 = nnTop_io_zout_1;
  assign T7 = nnTop_io_zout_0;
  assign io_yout = nnyout;
  assign T8 = T9;
  assign T9 = T11 + T10;
  assign T10 = nnTop_io_yout_11;
  assign T11 = T12;
  assign T12 = T13;
  assign T13 = T15 + T14;
  assign T14 = nnTop_io_yout_10;
  assign T15 = T16;
  assign T16 = T17;
  assign T17 = T19 + T18;
  assign T18 = nnTop_io_yout_9;
  assign T19 = T20;
  assign T20 = T21;
  assign T21 = T23 + T22;
  assign T22 = nnTop_io_yout_8;
  assign T23 = T24;
  assign T24 = T25;
  assign T25 = T27 + T26;
  assign T26 = nnTop_io_yout_7;
  assign T27 = T28;
  assign T28 = T29;
  assign T29 = T31 + T30;
  assign T30 = nnTop_io_yout_6;
  assign T31 = T32;
  assign T32 = T33;
  assign T33 = T35 + T34;
  assign T34 = nnTop_io_yout_5;
  assign T35 = T36;
  assign T36 = T37;
  assign T37 = T39 + T38;
  assign T38 = nnTop_io_yout_4;
  assign T39 = T40;
  assign T40 = T41;
  assign T41 = T43 + T42;
  assign T42 = nnTop_io_yout_3;
  assign T43 = T44;
  assign T44 = T45;
  assign T45 = T47 + T46;
  assign T46 = nnTop_io_yout_2;
  assign T47 = T48;
  assign T48 = T49;
  assign T49 = T51 + T50;
  assign T50 = nnTop_io_yout_1;
  assign T51 = nnTop_io_yout_0;
  assign io_xout = nnxout;
  assign T52 = T53;
  assign T53 = T55 + T54;
  assign T54 = nnTop_io_xout_2;
  assign T55 = T56;
  assign T56 = T57;
  assign T57 = T59 + T58;
  assign T58 = nnTop_io_xout_1;
  assign T59 = nnTop_io_xout_0;
  NN1Top nnTop(.clk(clk),
       .io_x_2( io_x ),
       .io_x_1( xShift_1 ),
       .io_x_0( xShift_0 ),
       .io_y_11( io_y ),
       .io_y_10( yShift_10 ),
       .io_y_9( yShift_9 ),
       .io_y_8( yShift_8 ),
       .io_y_7( yShift_7 ),
       .io_y_6( yShift_6 ),
       .io_y_5( yShift_5 ),
       .io_y_4( yShift_4 ),
       .io_y_3( yShift_3 ),
       .io_y_2( yShift_2 ),
       .io_y_1( yShift_1 ),
       .io_y_0( yShift_0 ),
       .io_z_2( io_z ),
       .io_z_1( zShift_1 ),
       .io_z_0( zShift_0 ),
       .io_b_11( io_b ),
       .io_b_10( bShift_10 ),
       .io_b_9( bShift_9 ),
       .io_b_8( bShift_8 ),
       .io_b_7( bShift_7 ),
       .io_b_6( bShift_6 ),
       .io_b_5( bShift_5 ),
       .io_b_4( bShift_4 ),
       .io_b_3( bShift_3 ),
       .io_b_2( bShift_2 ),
       .io_b_1( bShift_1 ),
       .io_b_0( bShift_0 ),
       .io_a_11_2( io_a ),
       .io_a_11_1( io_a ),
       .io_a_11_0( io_a ),
       .io_a_10_2( aShift_10_2 ),
       .io_a_10_1( aShift_10_1 ),
       .io_a_10_0( aShift_10_0 ),
       .io_a_9_2( aShift_9_2 ),
       .io_a_9_1( aShift_9_1 ),
       .io_a_9_0( aShift_9_0 ),
       .io_a_8_2( aShift_8_2 ),
       .io_a_8_1( aShift_8_1 ),
       .io_a_8_0( aShift_8_0 ),
       .io_a_7_2( aShift_7_2 ),
       .io_a_7_1( aShift_7_1 ),
       .io_a_7_0( aShift_7_0 ),
       .io_a_6_2( aShift_6_2 ),
       .io_a_6_1( aShift_6_1 ),
       .io_a_6_0( aShift_6_0 ),
       .io_a_5_2( aShift_5_2 ),
       .io_a_5_1( aShift_5_1 ),
       .io_a_5_0( aShift_5_0 ),
       .io_a_4_2( aShift_4_2 ),
       .io_a_4_1( aShift_4_1 ),
       .io_a_4_0( aShift_4_0 ),
       .io_a_3_2( aShift_3_2 ),
       .io_a_3_1( aShift_3_1 ),
       .io_a_3_0( aShift_3_0 ),
       .io_a_2_2( aShift_2_2 ),
       .io_a_2_1( aShift_2_1 ),
       .io_a_2_0( aShift_2_0 ),
       .io_a_1_2( aShift_1_2 ),
       .io_a_1_1( aShift_1_1 ),
       .io_a_1_0( aShift_1_0 ),
       .io_a_0_2( aShift_0_2 ),
       .io_a_0_1( aShift_0_1 ),
       .io_a_0_0( aShift_0_0 ),
       .io_c_2_2( io_c ),
       .io_c_2_1( io_c ),
       .io_c_2_0( io_c ),
       .io_c_1_2( cShift_1_2 ),
       .io_c_1_1( cShift_1_1 ),
       .io_c_1_0( cShift_1_0 ),
       .io_c_0_2( cShift_0_2 ),
       .io_c_0_1( cShift_0_1 ),
       .io_c_0_0( cShift_0_0 ),
       .io_lbda( io_lbda ),
       .io_xout_2( nnTop_io_xout_2 ),
       .io_xout_1( nnTop_io_xout_1 ),
       .io_xout_0( nnTop_io_xout_0 ),
       .io_yout_11( nnTop_io_yout_11 ),
       .io_yout_10( nnTop_io_yout_10 ),
       .io_yout_9( nnTop_io_yout_9 ),
       .io_yout_8( nnTop_io_yout_8 ),
       .io_yout_7( nnTop_io_yout_7 ),
       .io_yout_6( nnTop_io_yout_6 ),
       .io_yout_5( nnTop_io_yout_5 ),
       .io_yout_4( nnTop_io_yout_4 ),
       .io_yout_3( nnTop_io_yout_3 ),
       .io_yout_2( nnTop_io_yout_2 ),
       .io_yout_1( nnTop_io_yout_1 ),
       .io_yout_0( nnTop_io_yout_0 ),
       .io_zout_2( nnTop_io_zout_2 ),
       .io_zout_1( nnTop_io_zout_1 ),
       .io_zout_0( nnTop_io_zout_0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      cShift_0_0 <= 18'h0;
    end else begin
      cShift_0_0 <= cShift_1_0;
    end
    if(reset) begin
      cShift_1_0 <= 18'h0;
    end else begin
      cShift_1_0 <= cShift_2_0;
    end
    if(reset) begin
      cShift_2_0 <= 18'h0;
    end else begin
      cShift_2_0 <= io_c;
    end
    if(reset) begin
      cShift_0_1 <= 18'h0;
    end else begin
      cShift_0_1 <= cShift_1_1;
    end
    if(reset) begin
      cShift_1_1 <= 18'h0;
    end else begin
      cShift_1_1 <= cShift_2_1;
    end
    if(reset) begin
      cShift_2_1 <= 18'h0;
    end else begin
      cShift_2_1 <= io_c;
    end
    if(reset) begin
      cShift_0_2 <= 18'h0;
    end else begin
      cShift_0_2 <= cShift_1_2;
    end
    if(reset) begin
      cShift_1_2 <= 18'h0;
    end else begin
      cShift_1_2 <= cShift_2_2;
    end
    if(reset) begin
      cShift_2_2 <= 18'h0;
    end else begin
      cShift_2_2 <= io_c;
    end
    if(reset) begin
      aShift_0_0 <= 18'h0;
    end else begin
      aShift_0_0 <= aShift_1_0;
    end
    if(reset) begin
      aShift_1_0 <= 18'h0;
    end else begin
      aShift_1_0 <= aShift_2_0;
    end
    if(reset) begin
      aShift_2_0 <= 18'h0;
    end else begin
      aShift_2_0 <= aShift_3_0;
    end
    if(reset) begin
      aShift_3_0 <= 18'h0;
    end else begin
      aShift_3_0 <= aShift_4_0;
    end
    if(reset) begin
      aShift_4_0 <= 18'h0;
    end else begin
      aShift_4_0 <= aShift_5_0;
    end
    if(reset) begin
      aShift_5_0 <= 18'h0;
    end else begin
      aShift_5_0 <= aShift_6_0;
    end
    if(reset) begin
      aShift_6_0 <= 18'h0;
    end else begin
      aShift_6_0 <= aShift_7_0;
    end
    if(reset) begin
      aShift_7_0 <= 18'h0;
    end else begin
      aShift_7_0 <= aShift_8_0;
    end
    if(reset) begin
      aShift_8_0 <= 18'h0;
    end else begin
      aShift_8_0 <= aShift_9_0;
    end
    if(reset) begin
      aShift_9_0 <= 18'h0;
    end else begin
      aShift_9_0 <= aShift_10_0;
    end
    if(reset) begin
      aShift_10_0 <= 18'h0;
    end else begin
      aShift_10_0 <= aShift_11_0;
    end
    if(reset) begin
      aShift_11_0 <= 18'h0;
    end else begin
      aShift_11_0 <= io_a;
    end
    if(reset) begin
      aShift_0_1 <= 18'h0;
    end else begin
      aShift_0_1 <= aShift_1_1;
    end
    if(reset) begin
      aShift_1_1 <= 18'h0;
    end else begin
      aShift_1_1 <= aShift_2_1;
    end
    if(reset) begin
      aShift_2_1 <= 18'h0;
    end else begin
      aShift_2_1 <= aShift_3_1;
    end
    if(reset) begin
      aShift_3_1 <= 18'h0;
    end else begin
      aShift_3_1 <= aShift_4_1;
    end
    if(reset) begin
      aShift_4_1 <= 18'h0;
    end else begin
      aShift_4_1 <= aShift_5_1;
    end
    if(reset) begin
      aShift_5_1 <= 18'h0;
    end else begin
      aShift_5_1 <= aShift_6_1;
    end
    if(reset) begin
      aShift_6_1 <= 18'h0;
    end else begin
      aShift_6_1 <= aShift_7_1;
    end
    if(reset) begin
      aShift_7_1 <= 18'h0;
    end else begin
      aShift_7_1 <= aShift_8_1;
    end
    if(reset) begin
      aShift_8_1 <= 18'h0;
    end else begin
      aShift_8_1 <= aShift_9_1;
    end
    if(reset) begin
      aShift_9_1 <= 18'h0;
    end else begin
      aShift_9_1 <= aShift_10_1;
    end
    if(reset) begin
      aShift_10_1 <= 18'h0;
    end else begin
      aShift_10_1 <= aShift_11_1;
    end
    if(reset) begin
      aShift_11_1 <= 18'h0;
    end else begin
      aShift_11_1 <= io_a;
    end
    if(reset) begin
      aShift_0_2 <= 18'h0;
    end else begin
      aShift_0_2 <= aShift_1_2;
    end
    if(reset) begin
      aShift_1_2 <= 18'h0;
    end else begin
      aShift_1_2 <= aShift_2_2;
    end
    if(reset) begin
      aShift_2_2 <= 18'h0;
    end else begin
      aShift_2_2 <= aShift_3_2;
    end
    if(reset) begin
      aShift_3_2 <= 18'h0;
    end else begin
      aShift_3_2 <= aShift_4_2;
    end
    if(reset) begin
      aShift_4_2 <= 18'h0;
    end else begin
      aShift_4_2 <= aShift_5_2;
    end
    if(reset) begin
      aShift_5_2 <= 18'h0;
    end else begin
      aShift_5_2 <= aShift_6_2;
    end
    if(reset) begin
      aShift_6_2 <= 18'h0;
    end else begin
      aShift_6_2 <= aShift_7_2;
    end
    if(reset) begin
      aShift_7_2 <= 18'h0;
    end else begin
      aShift_7_2 <= aShift_8_2;
    end
    if(reset) begin
      aShift_8_2 <= 18'h0;
    end else begin
      aShift_8_2 <= aShift_9_2;
    end
    if(reset) begin
      aShift_9_2 <= 18'h0;
    end else begin
      aShift_9_2 <= aShift_10_2;
    end
    if(reset) begin
      aShift_10_2 <= 18'h0;
    end else begin
      aShift_10_2 <= aShift_11_2;
    end
    if(reset) begin
      aShift_11_2 <= 18'h0;
    end else begin
      aShift_11_2 <= io_a;
    end
    if(reset) begin
      bShift_0 <= 18'h0;
    end else begin
      bShift_0 <= bShift_1;
    end
    if(reset) begin
      bShift_1 <= 18'h0;
    end else begin
      bShift_1 <= bShift_2;
    end
    if(reset) begin
      bShift_2 <= 18'h0;
    end else begin
      bShift_2 <= bShift_3;
    end
    if(reset) begin
      bShift_3 <= 18'h0;
    end else begin
      bShift_3 <= bShift_4;
    end
    if(reset) begin
      bShift_4 <= 18'h0;
    end else begin
      bShift_4 <= bShift_5;
    end
    if(reset) begin
      bShift_5 <= 18'h0;
    end else begin
      bShift_5 <= bShift_6;
    end
    if(reset) begin
      bShift_6 <= 18'h0;
    end else begin
      bShift_6 <= bShift_7;
    end
    if(reset) begin
      bShift_7 <= 18'h0;
    end else begin
      bShift_7 <= bShift_8;
    end
    if(reset) begin
      bShift_8 <= 18'h0;
    end else begin
      bShift_8 <= bShift_9;
    end
    if(reset) begin
      bShift_9 <= 18'h0;
    end else begin
      bShift_9 <= bShift_10;
    end
    if(reset) begin
      bShift_10 <= 18'h0;
    end else begin
      bShift_10 <= bShift_11;
    end
    if(reset) begin
      bShift_11 <= 18'h0;
    end else begin
      bShift_11 <= io_b;
    end
    if(reset) begin
      zShift_0 <= 18'h0;
    end else begin
      zShift_0 <= zShift_1;
    end
    if(reset) begin
      zShift_1 <= 18'h0;
    end else begin
      zShift_1 <= zShift_2;
    end
    if(reset) begin
      zShift_2 <= 18'h0;
    end else begin
      zShift_2 <= io_z;
    end
    if(reset) begin
      yShift_0 <= 18'h0;
    end else begin
      yShift_0 <= yShift_1;
    end
    if(reset) begin
      yShift_1 <= 18'h0;
    end else begin
      yShift_1 <= yShift_2;
    end
    if(reset) begin
      yShift_2 <= 18'h0;
    end else begin
      yShift_2 <= yShift_3;
    end
    if(reset) begin
      yShift_3 <= 18'h0;
    end else begin
      yShift_3 <= yShift_4;
    end
    if(reset) begin
      yShift_4 <= 18'h0;
    end else begin
      yShift_4 <= yShift_5;
    end
    if(reset) begin
      yShift_5 <= 18'h0;
    end else begin
      yShift_5 <= yShift_6;
    end
    if(reset) begin
      yShift_6 <= 18'h0;
    end else begin
      yShift_6 <= yShift_7;
    end
    if(reset) begin
      yShift_7 <= 18'h0;
    end else begin
      yShift_7 <= yShift_8;
    end
    if(reset) begin
      yShift_8 <= 18'h0;
    end else begin
      yShift_8 <= yShift_9;
    end
    if(reset) begin
      yShift_9 <= 18'h0;
    end else begin
      yShift_9 <= yShift_10;
    end
    if(reset) begin
      yShift_10 <= 18'h0;
    end else begin
      yShift_10 <= yShift_11;
    end
    if(reset) begin
      yShift_11 <= 18'h0;
    end else begin
      yShift_11 <= io_y;
    end
    if(reset) begin
      xShift_0 <= 18'h0;
    end else begin
      xShift_0 <= xShift_1;
    end
    if(reset) begin
      xShift_1 <= 18'h0;
    end else begin
      xShift_1 <= xShift_2;
    end
    if(reset) begin
      xShift_2 <= 18'h0;
    end else begin
      xShift_2 <= io_x;
    end
    nnzout <= T0;
    nnyout <= T8;
    nnxout <= T52;
  end
endmodule

